sram_add_entry(0, 1, 0, 4, 128'h7ab000000000000000000deadbf);
sram_add_entry(0, 1, 4, 4, 128'h40200000000000000000093d46a);
sram_add_entry(0, 1, 8, 4, 128'h402000000000000000000d2356f);
sram_add_entry(0, 1, 12, 4, 128'h402000000000000000000676259);
sram_add_entry(0, 1, 16, 4, 128'h40200000000000000000046079b);
sram_add_entry(0, 1, 20, 4, 128'h4020000000000000000008c8892);
sram_add_entry(0, 1, 24, 4, 128'h40200000000000000000017cf44);
sram_add_entry(0, 1, 28, 4, 128'h402000000000000000000bc724b);
sram_add_entry(0, 1, 32, 4, 128'h402000000000000000000e97981);
sram_add_entry(0, 1, 36, 4, 128'h40200000000000000000077a9de);
sram_add_entry(0, 1, 40, 4, 128'h4020000000000000000002b7a6c);
sram_add_entry(0, 1, 44, 4, 128'h402000000000000000000504864);
sram_add_entry(0, 1, 48, 4, 128'h4020000000000000000008c6bb5);
sram_add_entry(0, 1, 52, 4, 128'h4020000000000000000007afada);
sram_add_entry(0, 1, 56, 4, 128'h402000000000000000000cc3650);
sram_add_entry(0, 1, 60, 4, 128'h40200000000000000000000dde1);
sram_add_entry(0, 1, 64, 4, 128'h40200000000000000000041bae2);
sram_add_entry(0, 1, 68, 4, 128'h4020000000000000000004b4f80);
sram_add_entry(0, 1, 72, 4, 128'h402000000000000000000ccad23);
sram_add_entry(0, 1, 76, 4, 128'h402000000000000000000987d18);
sram_add_entry(0, 1, 80, 4, 128'h402000000000000000000354214);
sram_add_entry(0, 1, 84, 4, 128'h4020000000000000000001b5bf0);
sram_add_entry(0, 1, 88, 4, 128'h402000000000000000000cfcfe0);
sram_add_entry(0, 1, 92, 4, 128'h4020000000000000000005dfdd7);
sram_add_entry(0, 1, 96, 4, 128'h402000000000000000000f65193);
sram_add_entry(0, 1, 100, 4, 128'h402000000000000000000699932);
sram_add_entry(0, 1, 104, 4, 128'h4020000000000000000003c1356);
sram_add_entry(0, 1, 108, 4, 128'h402000000000000000000da35e5);
sram_add_entry(0, 1, 112, 4, 128'h402000000000000000000ab08c2);
sram_add_entry(0, 1, 116, 4, 128'h40200000000000000000055162c);
sram_add_entry(0, 1, 120, 4, 128'h40200000000000000000048ac99);
sram_add_entry(0, 1, 124, 4, 128'h402000000000000000000cf2b64);
sram_add_entry(0, 1, 128, 4, 128'h402000000000000000000e09d8f);
sram_add_entry(0, 1, 132, 4, 128'h4020000000000000000001d11e0);
sram_add_entry(0, 1, 136, 4, 128'h402000000000000000000dc6d6f);
sram_add_entry(0, 1, 140, 4, 128'h40200000000000000000051d87e);
sram_add_entry(0, 1, 144, 4, 128'h402000000000000000000a23c19);
sram_add_entry(0, 1, 148, 4, 128'h402000000000000000000a8d569);
sram_add_entry(0, 1, 152, 4, 128'h4020000000000000000009d9ed7);
sram_add_entry(0, 1, 156, 4, 128'h40200000000000000000040e4d5);
sram_add_entry(0, 1, 160, 4, 128'h4020000000000000000006b550f);
sram_add_entry(0, 1, 164, 4, 128'h402000000000000000000b29e2e);
sram_add_entry(0, 1, 168, 4, 128'h4020000000000000000002e7cf1);
sram_add_entry(0, 1, 172, 4, 128'h4020000000000000000009200e3);
sram_add_entry(0, 1, 176, 4, 128'h402000000000000000000d9b933);
sram_add_entry(0, 1, 180, 4, 128'h402000000000000000000ed726f);
sram_add_entry(0, 1, 184, 4, 128'h4020000000000000000005a968d);
sram_add_entry(0, 1, 188, 4, 128'h402000000000000000000aa89df);
sram_add_entry(0, 1, 192, 4, 128'h402000000000000000000c1a0ac);
sram_add_entry(0, 1, 196, 4, 128'h402000000000000000000281727);
sram_add_entry(0, 1, 200, 4, 128'h402000000000000000000fe964b);
sram_add_entry(0, 1, 204, 4, 128'h402000000000000000000649d6a);
sram_add_entry(0, 1, 208, 4, 128'h402000000000000000000b66d0f);
sram_add_entry(0, 1, 212, 4, 128'h402000000000000000000a77176);
sram_add_entry(0, 1, 216, 4, 128'h402000000000000000000ab9e57);
sram_add_entry(0, 1, 220, 4, 128'h402000000000000000000e15190);
sram_add_entry(0, 1, 224, 4, 128'h402000000000000000000935b3f);
sram_add_entry(0, 1, 228, 4, 128'h40200000000000000000007d3e7);
sram_add_entry(0, 1, 232, 4, 128'h402000000000000000000d866b3);
sram_add_entry(0, 1, 236, 4, 128'h4020000000000000000004d2d96);
sram_add_entry(0, 1, 240, 4, 128'h402000000000000000000932137);
sram_add_entry(0, 1, 244, 4, 128'h402000000000000000000d76cda);
sram_add_entry(0, 1, 248, 4, 128'h402000000000000000000cfb810);
sram_add_entry(0, 1, 252, 4, 128'h4020000000000000000001f5e6f);
sram_add_entry(0, 1, 256, 4, 128'h4020000000000000000000866e5);
sram_add_entry(0, 1, 260, 4, 128'h402000000000000000000552409);
sram_add_entry(0, 1, 264, 4, 128'h40200000000000000000006819a);
sram_add_entry(0, 1, 268, 4, 128'h402000000000000000000dabaa8);
sram_add_entry(0, 1, 272, 4, 128'h4020000000000000000002fc8a9);
sram_add_entry(0, 1, 276, 4, 128'h4020000000000000000005014e0);
sram_add_entry(0, 1, 280, 4, 128'h402000000000000000000cc782f);
sram_add_entry(0, 1, 284, 4, 128'h4020000000000000000006dae2a);
sram_add_entry(0, 1, 288, 4, 128'h40200000000000000000039b496);
sram_add_entry(0, 1, 292, 4, 128'h4020000000000000000001cae91);
sram_add_entry(0, 1, 296, 4, 128'h402000000000000000000caff50);
sram_add_entry(0, 1, 300, 4, 128'h402000000000000000000033bd4);
sram_add_entry(0, 1, 304, 4, 128'h4020000000000000000004cb006);
sram_add_entry(0, 1, 308, 4, 128'h402000000000000000000a72599);
sram_add_entry(0, 1, 312, 4, 128'h40200000000000000000019efb1);
sram_add_entry(0, 1, 316, 4, 128'h402000000000000000000bc0688);
sram_add_entry(0, 1, 320, 4, 128'h40200000000000000000037cb96);
sram_add_entry(0, 1, 324, 4, 128'h40200000000000000000065d77e);
sram_add_entry(0, 1, 328, 4, 128'h402000000000000000000a4e182);
sram_add_entry(0, 1, 332, 4, 128'h402000000000000000000f9664b);
sram_add_entry(0, 1, 336, 4, 128'h402000000000000000000d9d504);
sram_add_entry(0, 1, 340, 4, 128'h402000000000000000000ac6429);
sram_add_entry(0, 1, 344, 4, 128'h4020000000000000000000587b1);
sram_add_entry(0, 1, 348, 4, 128'h40200000000000000000070b9ff);
sram_add_entry(0, 1, 352, 4, 128'h4020000000000000000007817b3);
sram_add_entry(0, 1, 356, 4, 128'h4020000000000000000005309c8);
sram_add_entry(0, 1, 360, 4, 128'h402000000000000000000263667);
sram_add_entry(0, 1, 364, 4, 128'h402000000000000000000baef4d);
sram_add_entry(0, 1, 368, 4, 128'h4020000000000000000009fe398);
sram_add_entry(0, 1, 372, 4, 128'h402000000000000000000f404b2);
sram_add_entry(0, 1, 376, 4, 128'h402000000000000000000e66811);
sram_add_entry(0, 1, 380, 4, 128'h4020000000000000000006c4854);
sram_add_entry(0, 1, 384, 4, 128'h402000000000000000000e41fbe);
sram_add_entry(0, 1, 388, 4, 128'h402000000000000000000ae926c);
sram_add_entry(0, 1, 392, 4, 128'h4020000000000000000008b4995);
sram_add_entry(0, 1, 396, 4, 128'h402000000000000000000ad9ee1);
sram_add_entry(0, 1, 400, 4, 128'h402000000000000000000e9cab6);
sram_add_entry(0, 1, 404, 4, 128'h402000000000000000000190690);
sram_add_entry(0, 1, 408, 4, 128'h402000000000000000000644cd1);
sram_add_entry(0, 1, 412, 4, 128'h402000000000000000000193143);
sram_add_entry(0, 1, 416, 4, 128'h402000000000000000000b38da9);
sram_add_entry(0, 1, 420, 4, 128'h402000000000000000000ad42fb);
sram_add_entry(0, 1, 424, 4, 128'h402000000000000000000f0c8e9);
sram_add_entry(0, 1, 428, 4, 128'h402000000000000000000c63e22);
sram_add_entry(0, 1, 432, 4, 128'h402000000000000000000ceae4f);
sram_add_entry(0, 1, 436, 4, 128'h40200000000000000000081fce1);
sram_add_entry(0, 1, 440, 4, 128'h4020000000000000000006c8b8a);
sram_add_entry(0, 1, 444, 4, 128'h402000000000000000000c9c607);
sram_add_entry(0, 1, 448, 4, 128'h40200000000000000000084f36d);
sram_add_entry(0, 1, 452, 4, 128'h402000000000000000000476c8a);
sram_add_entry(0, 1, 456, 4, 128'h402000000000000000000d0a28d);
sram_add_entry(0, 1, 460, 4, 128'h402000000000000000000a88374);
sram_add_entry(0, 1, 464, 4, 128'h402000000000000000000ec0149);
sram_add_entry(0, 1, 468, 4, 128'h402000000000000000000d54c20);
sram_add_entry(0, 1, 472, 4, 128'h402000000000000000000990140);
sram_add_entry(0, 1, 476, 4, 128'h402000000000000000000d8c32b);
sram_add_entry(0, 1, 480, 4, 128'h4020000000000000000009db7f1);
sram_add_entry(0, 1, 484, 4, 128'h4020000000000000000004fa872);
sram_add_entry(0, 1, 488, 4, 128'h402000000000000000000fa834c);
sram_add_entry(0, 1, 492, 4, 128'h402000000000000000000640129);
sram_add_entry(0, 1, 496, 4, 128'h402000000000000000000472ab0);
sram_add_entry(0, 1, 500, 4, 128'h402000000000000000000de8fce);
sram_add_entry(0, 1, 504, 4, 128'h402000000000000000000e5dd77);
sram_add_entry(0, 1, 508, 4, 128'h402000000000000000000e2e528);
sram_add_entry(0, 1, 512, 4, 128'h402000000000000000000c4a88f);
sram_add_entry(0, 1, 516, 4, 128'h40200000000000000000036d132);
sram_add_entry(0, 1, 520, 4, 128'h402000000000000000000103330);
sram_add_entry(0, 1, 524, 4, 128'h402000000000000000000210b4b);
sram_add_entry(0, 1, 528, 4, 128'h40200000000000000000023a29c);
sram_add_entry(0, 1, 532, 4, 128'h40200000000000000000018d134);
sram_add_entry(0, 1, 536, 4, 128'h402000000000000000000902d86);
sram_add_entry(0, 1, 540, 4, 128'h402000000000000000000599e1e);
sram_add_entry(0, 1, 544, 4, 128'h4020000000000000000008b80f3);
sram_add_entry(0, 1, 548, 4, 128'h402000000000000000000fdd6d9);
sram_add_entry(0, 1, 552, 4, 128'h402000000000000000000a822ed);
sram_add_entry(0, 1, 556, 4, 128'h402000000000000000000325c6b);
sram_add_entry(0, 1, 560, 4, 128'h402000000000000000000f3a0f1);
sram_add_entry(0, 1, 564, 4, 128'h40200000000000000000040625f);
sram_add_entry(0, 1, 568, 4, 128'h402000000000000000000062576);
sram_add_entry(0, 1, 572, 4, 128'h402000000000000000000247741);
sram_add_entry(0, 1, 576, 4, 128'h402000000000000000000e66076);
sram_add_entry(0, 1, 580, 4, 128'h402000000000000000000a1bfdb);
sram_add_entry(0, 1, 584, 4, 128'h402000000000000000000733a59);
sram_add_entry(0, 1, 588, 4, 128'h402000000000000000000d5364d);
sram_add_entry(0, 1, 592, 4, 128'h402000000000000000000bf32c7);
sram_add_entry(0, 1, 596, 4, 128'h402000000000000000000dc5dbf);
sram_add_entry(0, 1, 600, 4, 128'h4020000000000000000009a93fb);
sram_add_entry(0, 1, 604, 4, 128'h402000000000000000000cf1ba8);
sram_add_entry(0, 1, 608, 4, 128'h4020000000000000000002a29f0);
sram_add_entry(0, 1, 612, 4, 128'h402000000000000000000dbde8b);
sram_add_entry(0, 1, 616, 4, 128'h402000000000000000000009fe4);
sram_add_entry(0, 1, 620, 4, 128'h402000000000000000000180c0a);
sram_add_entry(0, 1, 624, 4, 128'h40200000000000000000088f835);
sram_add_entry(0, 1, 628, 4, 128'h40200000000000000000017109f);
sram_add_entry(0, 1, 632, 4, 128'h402000000000000000000889713);
sram_add_entry(0, 1, 636, 4, 128'h40200000000000000000041b6b6);
sram_add_entry(0, 1, 640, 4, 128'h402000000000000000000864de9);
sram_add_entry(0, 1, 644, 4, 128'h40200000000000000000007abce);
sram_add_entry(0, 1, 648, 4, 128'h402000000000000000000e12c35);
sram_add_entry(0, 1, 652, 4, 128'h402000000000000000000301447);
sram_add_entry(0, 1, 656, 4, 128'h402000000000000000000076b32);
sram_add_entry(0, 1, 660, 4, 128'h4020000000000000000004b21b3);
sram_add_entry(0, 1, 664, 4, 128'h402000000000000000000a87adb);
sram_add_entry(0, 1, 668, 4, 128'h4020000000000000000008e26bd);
sram_add_entry(0, 1, 672, 4, 128'h402000000000000000000e69464);
sram_add_entry(0, 1, 676, 4, 128'h402000000000000000000f1ae69);
sram_add_entry(0, 1, 680, 4, 128'h4020000000000000000003aec7a);
sram_add_entry(0, 1, 684, 4, 128'h402000000000000000000ee62e2);
sram_add_entry(0, 1, 688, 4, 128'h402000000000000000000e8bc68);
sram_add_entry(0, 1, 692, 4, 128'h4020000000000000000005b86a9);
sram_add_entry(0, 1, 696, 4, 128'h4020000000000000000007871a5);
sram_add_entry(0, 1, 700, 4, 128'h40200000000000000000055f1d9);
sram_add_entry(0, 1, 704, 4, 128'h40200000000000000000096e694);
sram_add_entry(0, 1, 708, 4, 128'h4020000000000000000001fe63b);
sram_add_entry(0, 1, 712, 4, 128'h402000000000000000000806547);
sram_add_entry(0, 1, 716, 4, 128'h40200000000000000000025c72f);
sram_add_entry(0, 1, 720, 4, 128'h402000000000000000000a62af6);
sram_add_entry(0, 1, 724, 4, 128'h4020000000000000000009d5417);
sram_add_entry(0, 1, 728, 4, 128'h4020000000000000000002c51af);
sram_add_entry(0, 1, 732, 4, 128'h4020000000000000000002f7ca4);
sram_add_entry(0, 1, 736, 4, 128'h402000000000000000000c3d2cf);
sram_add_entry(0, 1, 740, 4, 128'h4020000000000000000002f8d88);
sram_add_entry(0, 1, 744, 4, 128'h402000000000000000000128302);
sram_add_entry(0, 1, 748, 4, 128'h4020000000000000000003cc6e7);
sram_add_entry(0, 1, 752, 4, 128'h402000000000000000000bebdfb);
sram_add_entry(0, 1, 756, 4, 128'h402000000000000000000aaacbb);
sram_add_entry(0, 1, 760, 4, 128'h40200000000000000000035afca);
sram_add_entry(0, 1, 764, 4, 128'h4020000000000000000003f635d);
sram_add_entry(0, 1, 768, 4, 128'h4020000000000000000009dc27f);
sram_add_entry(0, 1, 772, 4, 128'h402000000000000000000f64438);
sram_add_entry(0, 1, 776, 4, 128'h4020000000000000000001cde19);
sram_add_entry(0, 1, 780, 4, 128'h402000000000000000000ad0b70);
sram_add_entry(0, 1, 784, 4, 128'h402000000000000000000b2a22c);
sram_add_entry(0, 1, 788, 4, 128'h402000000000000000000c40815);
sram_add_entry(0, 1, 792, 4, 128'h402000000000000000000a08a15);
sram_add_entry(0, 1, 796, 4, 128'h402000000000000000000294352);
sram_add_entry(0, 1, 800, 4, 128'h40200000000000000000009f922);
sram_add_entry(0, 1, 804, 4, 128'h402000000000000000000c44933);
sram_add_entry(0, 1, 808, 4, 128'h402000000000000000000cba9fb);
sram_add_entry(0, 1, 812, 4, 128'h402000000000000000000cee397);
sram_add_entry(0, 1, 816, 4, 128'h4020000000000000000005ab855);
sram_add_entry(0, 1, 820, 4, 128'h402000000000000000000c37cff);
sram_add_entry(0, 1, 824, 4, 128'h4020000000000000000000f1815);
sram_add_entry(0, 1, 828, 4, 128'h4020000000000000000001fecf8);
sram_add_entry(0, 1, 832, 4, 128'h4020000000000000000002f0cd3);
sram_add_entry(0, 1, 836, 4, 128'h402000000000000000000cdfdc7);
sram_add_entry(0, 1, 840, 4, 128'h402000000000000000000eada3f);
sram_add_entry(0, 1, 844, 4, 128'h402000000000000000000c5239f);
sram_add_entry(0, 1, 848, 4, 128'h4020000000000000000002e0306);
sram_add_entry(0, 1, 852, 4, 128'h4020000000000000000009b50e8);
sram_add_entry(0, 1, 856, 4, 128'h402000000000000000000244d2d);
sram_add_entry(0, 1, 860, 4, 128'h402000000000000000000d04cf1);
sram_add_entry(0, 1, 864, 4, 128'h40200000000000000000012056a);
sram_add_entry(0, 1, 868, 4, 128'h40200000000000000000017ca62);
sram_add_entry(0, 1, 872, 4, 128'h4020000000000000000003f7a75);
sram_add_entry(0, 1, 876, 4, 128'h4020000000000000000007a839f);
sram_add_entry(0, 1, 880, 4, 128'h4020000000000000000000488d5);
sram_add_entry(0, 1, 884, 4, 128'h40200000000000000000034ae81);
sram_add_entry(0, 1, 888, 4, 128'h4020000000000000000001ee202);
sram_add_entry(0, 1, 892, 4, 128'h402000000000000000000183ea5);
sram_add_entry(0, 1, 896, 4, 128'h402000000000000000000c5cf43);
sram_add_entry(0, 1, 900, 4, 128'h402000000000000000000e2bc13);
sram_add_entry(0, 1, 904, 4, 128'h4020000000000000000001fd051);
sram_add_entry(0, 1, 908, 4, 128'h4020000000000000000001d970f);
sram_add_entry(0, 1, 912, 4, 128'h402000000000000000000c403c7);
sram_add_entry(0, 1, 916, 4, 128'h40200000000000000000088f8af);
sram_add_entry(0, 1, 920, 4, 128'h402000000000000000000522f39);
sram_add_entry(0, 1, 924, 4, 128'h402000000000000000000f385d1);
sram_add_entry(0, 1, 928, 4, 128'h4020000000000000000009777c8);
sram_add_entry(0, 1, 932, 4, 128'h402000000000000000000ffee98);
sram_add_entry(0, 1, 936, 4, 128'h4020000000000000000008f8852);
sram_add_entry(0, 1, 940, 4, 128'h40200000000000000000022a823);
sram_add_entry(0, 1, 944, 4, 128'h402000000000000000000aabbdd);
sram_add_entry(0, 1, 948, 4, 128'h402000000000000000000c4d792);
sram_add_entry(0, 1, 952, 4, 128'h4020000000000000000001af82d);
sram_add_entry(0, 1, 956, 4, 128'h40200000000000000000012e62a);
sram_add_entry(0, 1, 960, 4, 128'h40200000000000000000084feb8);
sram_add_entry(0, 1, 964, 4, 128'h402000000000000000000e90935);
sram_add_entry(0, 1, 968, 4, 128'h402000000000000000000daeacf);
sram_add_entry(0, 1, 972, 4, 128'h402000000000000000000f7fb36);
sram_add_entry(0, 1, 976, 4, 128'h4020000000000000000000b754c);
sram_add_entry(0, 1, 980, 4, 128'h40200000000000000000072a0d2);
sram_add_entry(0, 1, 984, 4, 128'h40200000000000000000014c7a8);
sram_add_entry(0, 1, 988, 4, 128'h4020000000000000000002e7ccb);
sram_add_entry(0, 1, 992, 4, 128'h402000000000000000000172d6b);
sram_add_entry(0, 1, 996, 4, 128'h4020000000000000000005cbd69);
sram_add_entry(0, 1, 1000, 4, 128'h402000000000000000000838848);
sram_add_entry(0, 1, 1004, 4, 128'h402000000000000000000e57f48);
sram_add_entry(0, 1, 1008, 4, 128'h402000000000000000000879954);
sram_add_entry(0, 1, 1012, 4, 128'h4020000000000000000003f3b48);
sram_add_entry(0, 1, 1016, 4, 128'h402000000000000000000aa15a1);
sram_add_entry(0, 1, 1020, 4, 128'h40200000000000000000072e889);
sram_add_entry(0, 1, 1024, 4, 128'h40200000000000000000001b542);
sram_add_entry(0, 1, 1028, 4, 128'h402000000000000000000296632);
sram_add_entry(0, 1, 1032, 4, 128'h40200000000000000000038ad9e);
sram_add_entry(0, 1, 1036, 4, 128'h402000000000000000000dd5b20);
sram_add_entry(0, 1, 1040, 4, 128'h4020000000000000000007e3d3f);
sram_add_entry(0, 1, 1044, 4, 128'h402000000000000000000de577e);
sram_add_entry(0, 1, 1048, 4, 128'h4020000000000000000005f90c0);
sram_add_entry(0, 1, 1052, 4, 128'h402000000000000000000d30cb2);
sram_add_entry(0, 1, 1056, 4, 128'h4020000000000000000008ebe76);
sram_add_entry(0, 1, 1060, 4, 128'h4020000000000000000002d1e33);
sram_add_entry(0, 1, 1064, 4, 128'h40200000000000000000078e2fd);
sram_add_entry(0, 1, 1068, 4, 128'h4020000000000000000008595a0);
sram_add_entry(0, 1, 1072, 4, 128'h4020000000000000000004d7b60);
sram_add_entry(0, 1, 1076, 4, 128'h4020000000000000000000a5d4d);
sram_add_entry(0, 1, 1080, 4, 128'h402000000000000000000b6a7b0);
sram_add_entry(0, 1, 1084, 4, 128'h402000000000000000000b9d0d8);
sram_add_entry(0, 1, 1088, 4, 128'h4020000000000000000007c54d0);
sram_add_entry(0, 1, 1092, 4, 128'h402000000000000000000000fab);
sram_add_entry(0, 1, 1096, 4, 128'h402000000000000000000526452);
sram_add_entry(0, 1, 1100, 4, 128'h402000000000000000000eea715);
sram_add_entry(0, 1, 1104, 4, 128'h402000000000000000000b958bc);
sram_add_entry(0, 1, 1108, 4, 128'h402000000000000000000a9b50c);
sram_add_entry(0, 1, 1112, 4, 128'h402000000000000000000fcbf5c);
sram_add_entry(0, 1, 1116, 4, 128'h402000000000000000000d7128e);
sram_add_entry(0, 1, 1120, 4, 128'h402000000000000000000287b14);
sram_add_entry(0, 1, 1124, 4, 128'h40200000000000000000099d893);
sram_add_entry(0, 1, 1128, 4, 128'h402000000000000000000ce1be7);
sram_add_entry(0, 1, 1132, 4, 128'h402000000000000000000275c14);
sram_add_entry(0, 1, 1136, 4, 128'h402000000000000000000b2ecf6);
sram_add_entry(0, 1, 1140, 4, 128'h40200000000000000000032209f);
sram_add_entry(0, 1, 1144, 4, 128'h4020000000000000000008890e9);
sram_add_entry(0, 1, 1148, 4, 128'h4020000000000000000005df3a2);
sram_add_entry(0, 1, 1152, 4, 128'h402000000000000000000681f7e);
sram_add_entry(0, 1, 1156, 4, 128'h40200000000000000000052ac42);
sram_add_entry(0, 1, 1160, 4, 128'h40200000000000000000062b76d);
sram_add_entry(0, 1, 1164, 4, 128'h4020000000000000000002a3054);
sram_add_entry(0, 1, 1168, 4, 128'h402000000000000000000a6aacb);
sram_add_entry(0, 1, 1172, 4, 128'h402000000000000000000fad7b0);
sram_add_entry(0, 1, 1176, 4, 128'h402000000000000000000e45af7);
sram_add_entry(0, 1, 1180, 4, 128'h4020000000000000000001b8312);
sram_add_entry(0, 1, 1184, 4, 128'h4020000000000000000004d7686);
sram_add_entry(0, 1, 1188, 4, 128'h4020000000000000000009e9f11);
sram_add_entry(0, 1, 1192, 4, 128'h4020000000000000000003752b8);
sram_add_entry(0, 1, 1196, 4, 128'h4020000000000000000009fff19);
sram_add_entry(0, 1, 1200, 4, 128'h4020000000000000000003deeb0);
sram_add_entry(0, 1, 1204, 4, 128'h4020000000000000000004d0cc0);
sram_add_entry(0, 1, 1208, 4, 128'h402000000000000000000ad4e0b);
sram_add_entry(0, 1, 1212, 4, 128'h402000000000000000000d93c76);
sram_add_entry(0, 1, 1216, 4, 128'h402000000000000000000a363f3);
sram_add_entry(0, 1, 1220, 4, 128'h402000000000000000000fe7a4a);
sram_add_entry(0, 1, 1224, 4, 128'h4020000000000000000006750fd);
sram_add_entry(0, 1, 1228, 4, 128'h402000000000000000000fa4199);
sram_add_entry(0, 1, 1232, 4, 128'h402000000000000000000d91f85);
sram_add_entry(0, 1, 1236, 4, 128'h4020000000000000000006021c5);
sram_add_entry(0, 1, 1240, 4, 128'h402000000000000000000b7fc65);
sram_add_entry(0, 1, 1244, 4, 128'h4020000000000000000000d6e41);
sram_add_entry(0, 1, 1248, 4, 128'h4020000000000000000001fc6a1);
sram_add_entry(0, 1, 1252, 4, 128'h402000000000000000000d152b0);
sram_add_entry(0, 1, 1256, 4, 128'h4020000000000000000002f8780);
sram_add_entry(0, 1, 1260, 4, 128'h4020000000000000000000a9948);
sram_add_entry(0, 1, 1264, 4, 128'h402000000000000000000249ab8);
sram_add_entry(0, 1, 1268, 4, 128'h402000000000000000000472875);
sram_add_entry(0, 1, 1272, 4, 128'h4020000000000000000006d2196);
sram_add_entry(0, 1, 1276, 4, 128'h40200000000000000000010373f);
sram_add_entry(0, 1, 1280, 4, 128'h402000000000000000000c0f50e);
sram_add_entry(0, 1, 1284, 4, 128'h402000000000000000000dd84a8);
sram_add_entry(0, 1, 1288, 4, 128'h402000000000000000000324444);
sram_add_entry(0, 1, 1292, 4, 128'h402000000000000000000b11fe3);
sram_add_entry(0, 1, 1296, 4, 128'h402000000000000000000d3c003);
sram_add_entry(0, 1, 1300, 4, 128'h40200000000000000000022c068);
sram_add_entry(0, 1, 1304, 4, 128'h402000000000000000000200557);
sram_add_entry(0, 1, 1308, 4, 128'h402000000000000000000d760d5);
sram_add_entry(0, 1, 1312, 4, 128'h402000000000000000000404d84);
sram_add_entry(0, 1, 1316, 4, 128'h40200000000000000000038a6a0);
sram_add_entry(0, 1, 1320, 4, 128'h4020000000000000000003a4640);
sram_add_entry(0, 1, 1324, 4, 128'h4020000000000000000004a10b1);
sram_add_entry(0, 1, 1328, 4, 128'h402000000000000000000b30115);
sram_add_entry(0, 1, 1332, 4, 128'h4020000000000000000008aeaa5);
sram_add_entry(0, 1, 1336, 4, 128'h402000000000000000000f1cc59);
sram_add_entry(0, 1, 1340, 4, 128'h4020000000000000000007f6f35);
sram_add_entry(0, 1, 1344, 4, 128'h402000000000000000000465838);
sram_add_entry(0, 1, 1348, 4, 128'h402000000000000000000c08db5);
sram_add_entry(0, 1, 1352, 4, 128'h402000000000000000000fd7be1);
sram_add_entry(0, 1, 1356, 4, 128'h40200000000000000000000a0f3);
sram_add_entry(0, 1, 1360, 4, 128'h402000000000000000000b91869);
sram_add_entry(0, 1, 1364, 4, 128'h402000000000000000000c0ad63);
sram_add_entry(0, 1, 1368, 4, 128'h402000000000000000000b08e22);
sram_add_entry(0, 1, 1372, 4, 128'h402000000000000000000f68553);
sram_add_entry(0, 1, 1376, 4, 128'h40200000000000000000064927f);
sram_add_entry(0, 1, 1380, 4, 128'h40200000000000000000083a02e);
sram_add_entry(0, 1, 1384, 4, 128'h402000000000000000000be5a96);
sram_add_entry(0, 1, 1388, 4, 128'h4020000000000000000006e40d1);
sram_add_entry(0, 1, 1392, 4, 128'h402000000000000000000f76daa);
sram_add_entry(0, 1, 1396, 4, 128'h402000000000000000000260806);
sram_add_entry(0, 1, 1400, 4, 128'h402000000000000000000aaf348);
sram_add_entry(0, 1, 1404, 4, 128'h4020000000000000000000be1a7);
sram_add_entry(0, 1, 1408, 4, 128'h402000000000000000000a59283);
sram_add_entry(0, 1, 1412, 4, 128'h4020000000000000000009fd1ab);
sram_add_entry(0, 1, 1416, 4, 128'h4020000000000000000008acbff);
sram_add_entry(0, 1, 1420, 4, 128'h4020000000000000000004deca7);
sram_add_entry(0, 1, 1424, 4, 128'h40200000000000000000028e13a);
sram_add_entry(0, 1, 1428, 4, 128'h402000000000000000000a299ca);
sram_add_entry(0, 1, 1432, 4, 128'h40200000000000000000099a477);
sram_add_entry(0, 1, 1436, 4, 128'h40200000000000000000044a766);
sram_add_entry(0, 1, 1440, 4, 128'h402000000000000000000d3a394);
sram_add_entry(0, 1, 1444, 4, 128'h402000000000000000000ecc3e8);
sram_add_entry(0, 1, 1448, 4, 128'h402000000000000000000ebab0e);
sram_add_entry(0, 1, 1452, 4, 128'h4020000000000000000007f07a0);
sram_add_entry(0, 1, 1456, 4, 128'h4020000000000000000001940da);
sram_add_entry(0, 1, 1460, 4, 128'h402000000000000000000dd77fd);
sram_add_entry(0, 1, 1464, 4, 128'h40200000000000000000027a422);
sram_add_entry(0, 1, 1468, 4, 128'h402000000000000000000e19559);
sram_add_entry(0, 1, 1472, 4, 128'h402000000000000000000008d63);
sram_add_entry(0, 1, 1476, 4, 128'h40200000000000000000001193c);
sram_add_entry(0, 1, 1480, 4, 128'h40200000000000000000046a7c0);
sram_add_entry(0, 1, 1484, 4, 128'h402000000000000000000c71745);
sram_add_entry(0, 1, 1488, 4, 128'h402000000000000000000ee0321);
sram_add_entry(0, 1, 1492, 4, 128'h40200000000000000000021c943);
sram_add_entry(0, 1, 1496, 4, 128'h4020000000000000000005334c6);
sram_add_entry(0, 1, 1500, 4, 128'h402000000000000000000cbd414);
sram_add_entry(0, 1, 1504, 4, 128'h402000000000000000000ab0538);
sram_add_entry(0, 1, 1508, 4, 128'h402000000000000000000f176c0);
sram_add_entry(0, 1, 1512, 4, 128'h4020000000000000000008512ed);
sram_add_entry(0, 1, 1516, 4, 128'h402000000000000000000a0128d);
sram_add_entry(0, 1, 1520, 4, 128'h402000000000000000000db3124);
sram_add_entry(0, 1, 1524, 4, 128'h4020000000000000000003d7888);
sram_add_entry(0, 1, 1528, 4, 128'h40200000000000000000006f91b);
sram_add_entry(0, 1, 1532, 4, 128'h402000000000000000000b21e43);
sram_add_entry(0, 1, 1536, 4, 128'h4020000000000000000008de00c);
sram_add_entry(0, 1, 1540, 4, 128'h402000000000000000000ad6a91);
sram_add_entry(0, 1, 1544, 4, 128'h4020000000000000000009982b5);
sram_add_entry(0, 1, 1548, 4, 128'h402000000000000000000f936b6);
sram_add_entry(0, 1, 1552, 4, 128'h402000000000000000000fb8434);
sram_add_entry(0, 1, 1556, 4, 128'h40200000000000000000061ac31);
sram_add_entry(0, 1, 1560, 4, 128'h402000000000000000000000d66);
sram_add_entry(0, 1, 1564, 4, 128'h402000000000000000000cb4d6b);
sram_add_entry(0, 1, 1568, 4, 128'h402000000000000000000952555);
sram_add_entry(0, 1, 1572, 4, 128'h402000000000000000000d662de);
sram_add_entry(0, 1, 1576, 4, 128'h402000000000000000000aa0ea6);
sram_add_entry(0, 1, 1580, 4, 128'h402000000000000000000ba2e0f);
sram_add_entry(0, 1, 1584, 4, 128'h402000000000000000000f7491c);
sram_add_entry(0, 1, 1588, 4, 128'h4020000000000000000008d68ee);
sram_add_entry(0, 1, 1592, 4, 128'h402000000000000000000a366a5);
sram_add_entry(0, 1, 1596, 4, 128'h4020000000000000000007672fe);
sram_add_entry(0, 1, 1600, 4, 128'h4020000000000000000004e0e5b);
sram_add_entry(0, 1, 1604, 4, 128'h402000000000000000000f69f93);
sram_add_entry(0, 1, 1608, 4, 128'h402000000000000000000dc64a3);
sram_add_entry(0, 1, 1612, 4, 128'h4020000000000000000003e36d7);
sram_add_entry(0, 1, 1616, 4, 128'h40200000000000000000020cd14);
sram_add_entry(0, 1, 1620, 4, 128'h402000000000000000000fd80ee);
sram_add_entry(0, 1, 1624, 4, 128'h40200000000000000000014a853);
sram_add_entry(0, 1, 1628, 4, 128'h402000000000000000000d34e71);
sram_add_entry(0, 1, 1632, 4, 128'h4020000000000000000004da43e);
sram_add_entry(0, 1, 1636, 4, 128'h4020000000000000000002dcdd0);
sram_add_entry(0, 1, 1640, 4, 128'h402000000000000000000ff51e4);
sram_add_entry(0, 1, 1644, 4, 128'h4020000000000000000005e4c3b);
sram_add_entry(0, 1, 1648, 4, 128'h402000000000000000000919a50);
sram_add_entry(0, 1, 1652, 4, 128'h40200000000000000000005c6f6);
sram_add_entry(0, 1, 1656, 4, 128'h4020000000000000000004880e1);
sram_add_entry(0, 1, 1660, 4, 128'h402000000000000000000b52f6e);
sram_add_entry(0, 1, 1664, 4, 128'h4020000000000000000006330f5);
sram_add_entry(0, 1, 1668, 4, 128'h40200000000000000000087589c);
sram_add_entry(0, 1, 1672, 4, 128'h402000000000000000000ae87c5);
sram_add_entry(0, 1, 1676, 4, 128'h40200000000000000000088b591);
sram_add_entry(0, 1, 1680, 4, 128'h402000000000000000000a9681c);
sram_add_entry(0, 1, 1684, 4, 128'h4020000000000000000005bfe8c);
sram_add_entry(0, 1, 1688, 4, 128'h402000000000000000000feeabb);
sram_add_entry(0, 1, 1692, 4, 128'h4020000000000000000005bfef3);
sram_add_entry(0, 1, 1696, 4, 128'h402000000000000000000c439f5);
sram_add_entry(0, 1, 1700, 4, 128'h402000000000000000000cbb611);
sram_add_entry(0, 1, 1704, 4, 128'h4020000000000000000006bf841);
sram_add_entry(0, 1, 1708, 4, 128'h40200000000000000000014eb96);
sram_add_entry(0, 1, 1712, 4, 128'h402000000000000000000cb6ce3);
sram_add_entry(0, 1, 1716, 4, 128'h402000000000000000000be0907);
sram_add_entry(0, 1, 1720, 4, 128'h402000000000000000000f515b5);
sram_add_entry(0, 1, 1724, 4, 128'h402000000000000000000d4b21b);
sram_add_entry(0, 1, 1728, 4, 128'h402000000000000000000aed1b5);
sram_add_entry(0, 1, 1732, 4, 128'h4020000000000000000000187e1);
sram_add_entry(0, 1, 1736, 4, 128'h4020000000000000000003bf896);
sram_add_entry(0, 1, 1740, 4, 128'h402000000000000000000d53055);
sram_add_entry(0, 1, 1744, 4, 128'h402000000000000000000d85a46);
sram_add_entry(0, 1, 1748, 4, 128'h402000000000000000000b70da5);
sram_add_entry(0, 1, 1752, 4, 128'h402000000000000000000f14efb);
sram_add_entry(0, 1, 1756, 4, 128'h402000000000000000000ceed54);
sram_add_entry(0, 1, 1760, 4, 128'h4020000000000000000001c63cc);
sram_add_entry(0, 1, 1764, 4, 128'h4020000000000000000002e657b);
sram_add_entry(0, 1, 1768, 4, 128'h4020000000000000000001b7bb1);
sram_add_entry(0, 1, 1772, 4, 128'h402000000000000000000a490bb);
sram_add_entry(0, 1, 1776, 4, 128'h40200000000000000000077f7c3);
sram_add_entry(0, 1, 1780, 4, 128'h402000000000000000000ce3879);
sram_add_entry(0, 1, 1784, 4, 128'h4020000000000000000003d62f7);
sram_add_entry(0, 1, 1788, 4, 128'h402000000000000000000d3c317);
sram_add_entry(0, 1, 1792, 4, 128'h402000000000000000000cd4052);
sram_add_entry(0, 1, 1796, 4, 128'h402000000000000000000366029);
sram_add_entry(0, 1, 1800, 4, 128'h402000000000000000000249c31);
sram_add_entry(0, 1, 1804, 4, 128'h402000000000000000000f85353);
sram_add_entry(0, 1, 1808, 4, 128'h402000000000000000000ba861d);
sram_add_entry(0, 1, 1812, 4, 128'h4020000000000000000007b4f14);
sram_add_entry(0, 1, 1816, 4, 128'h402000000000000000000e9a8b0);
sram_add_entry(0, 1, 1820, 4, 128'h40200000000000000000048daff);
sram_add_entry(0, 1, 1824, 4, 128'h40200000000000000000009eeb3);
sram_add_entry(0, 1, 1828, 4, 128'h40200000000000000000001ea67);
sram_add_entry(0, 1, 1832, 4, 128'h402000000000000000000b2c532);
sram_add_entry(0, 1, 1836, 4, 128'h4020000000000000000008cdabd);
sram_add_entry(0, 1, 1840, 4, 128'h402000000000000000000e33611);
sram_add_entry(0, 1, 1844, 4, 128'h402000000000000000000888646);
sram_add_entry(0, 1, 1848, 4, 128'h4020000000000000000007532ec);
sram_add_entry(0, 1, 1852, 4, 128'h402000000000000000000ef77eb);
sram_add_entry(0, 1, 1856, 4, 128'h402000000000000000000836a74);
sram_add_entry(0, 1, 1860, 4, 128'h40200000000000000000060abde);
sram_add_entry(0, 1, 1864, 4, 128'h4020000000000000000001fb207);
sram_add_entry(0, 1, 1868, 4, 128'h4020000000000000000001fd4bb);
sram_add_entry(0, 1, 1872, 4, 128'h402000000000000000000e37673);
sram_add_entry(0, 1, 1876, 4, 128'h402000000000000000000e78f3e);
sram_add_entry(0, 1, 1880, 4, 128'h402000000000000000000f089bc);
sram_add_entry(0, 1, 1884, 4, 128'h402000000000000000000989a46);
sram_add_entry(0, 1, 1888, 4, 128'h40200000000000000000004872d);
sram_add_entry(0, 1, 1892, 4, 128'h4020000000000000000007d4a59);
sram_add_entry(0, 1, 1896, 4, 128'h40200000000000000000079148c);
sram_add_entry(0, 1, 1900, 4, 128'h402000000000000000000ca4d53);
sram_add_entry(0, 1, 1904, 4, 128'h402000000000000000000318859);
sram_add_entry(0, 1, 1908, 4, 128'h402000000000000000000d19af7);
sram_add_entry(0, 1, 1912, 4, 128'h402000000000000000000270545);
sram_add_entry(0, 1, 1916, 4, 128'h40200000000000000000094a8f5);
sram_add_entry(0, 1, 1920, 4, 128'h402000000000000000000fd4a65);
sram_add_entry(0, 1, 1924, 4, 128'h40200000000000000000014a4ed);
sram_add_entry(0, 1, 1928, 4, 128'h402000000000000000000b279ba);
sram_add_entry(0, 1, 1932, 4, 128'h40200000000000000000063905b);
sram_add_entry(0, 1, 1936, 4, 128'h402000000000000000000528285);
sram_add_entry(0, 1, 1940, 4, 128'h402000000000000000000bd6eb1);
sram_add_entry(0, 1, 1944, 4, 128'h402000000000000000000136e6c);
sram_add_entry(0, 1, 1948, 4, 128'h4020000000000000000009b3456);
sram_add_entry(0, 1, 1952, 4, 128'h402000000000000000000254c0a);
sram_add_entry(0, 1, 1956, 4, 128'h402000000000000000000ec438c);
sram_add_entry(0, 1, 1960, 4, 128'h40200000000000000000084699d);
sram_add_entry(0, 1, 1964, 4, 128'h4020000000000000000000d0224);
sram_add_entry(0, 1, 1968, 4, 128'h402000000000000000000c49916);
sram_add_entry(0, 1, 1972, 4, 128'h402000000000000000000ff4173);
sram_add_entry(0, 1, 1976, 4, 128'h40200000000000000000081bccf);
sram_add_entry(0, 1, 1980, 4, 128'h4020000000000000000006fed17);
sram_add_entry(0, 1, 1984, 4, 128'h4020000000000000000002329d9);
sram_add_entry(0, 1, 1988, 4, 128'h402000000000000000000e35295);
sram_add_entry(0, 1, 1992, 4, 128'h40200000000000000000097a6ce);
sram_add_entry(0, 1, 1996, 4, 128'h4020000000000000000007355fd);
sram_add_entry(0, 1, 2000, 4, 128'h402000000000000000000b5e794);
sram_add_entry(0, 1, 2004, 4, 128'h4020000000000000000003295ab);
sram_add_entry(0, 1, 2008, 4, 128'h402000000000000000000eca5ce);
sram_add_entry(0, 1, 2012, 4, 128'h40200000000000000000087bf14);
sram_add_entry(0, 1, 2016, 4, 128'h402000000000000000000a166f5);
sram_add_entry(0, 1, 2020, 4, 128'h402000000000000000000c0b98a);
sram_add_entry(0, 1, 2024, 4, 128'h402000000000000000000452cdc);
sram_add_entry(0, 1, 2028, 4, 128'h40200000000000000000078e1e0);
sram_add_entry(0, 1, 2032, 4, 128'h40200000000000000000092eb8c);
sram_add_entry(0, 1, 2036, 4, 128'h402000000000000000000129629);
sram_add_entry(0, 1, 2040, 4, 128'h402000000000000000000bc837b);
sram_add_entry(0, 1, 2044, 4, 128'h4020000000000000000009cda8f);
sram_add_entry(0, 1, 2048, 4, 128'h4020000000000000000003e36f7);
sram_add_entry(0, 1, 2052, 4, 128'h4020000000000000000008a27cd);
sram_add_entry(0, 1, 2056, 4, 128'h402000000000000000000462c62);
sram_add_entry(0, 1, 2060, 4, 128'h402000000000000000000dfcade);
sram_add_entry(0, 1, 2064, 4, 128'h4020000000000000000008989c8);
sram_add_entry(0, 1, 2068, 4, 128'h4020000000000000000006c0294);
sram_add_entry(0, 1, 2072, 4, 128'h402000000000000000000bcd2eb);
sram_add_entry(0, 1, 2076, 4, 128'h4020000000000000000003bff68);
sram_add_entry(0, 1, 2080, 4, 128'h4020000000000000000006b9b27);
sram_add_entry(0, 1, 2084, 4, 128'h40200000000000000000022b3ea);
sram_add_entry(0, 1, 2088, 4, 128'h40200000000000000000041688a);
sram_add_entry(0, 1, 2092, 4, 128'h402000000000000000000e21345);
sram_add_entry(0, 1, 2096, 4, 128'h40200000000000000000073d32b);
sram_add_entry(0, 1, 2100, 4, 128'h402000000000000000000a2a953);
sram_add_entry(0, 1, 2104, 4, 128'h4020000000000000000004e430c);
sram_add_entry(0, 1, 2108, 4, 128'h40200000000000000000064d84c);
sram_add_entry(0, 1, 2112, 4, 128'h4020000000000000000002f0b4c);
sram_add_entry(0, 1, 2116, 4, 128'h4020000000000000000003b69f1);
sram_add_entry(0, 1, 2120, 4, 128'h4020000000000000000000ac0c0);
sram_add_entry(0, 1, 2124, 4, 128'h40200000000000000000002cb8c);
sram_add_entry(0, 1, 2128, 4, 128'h402000000000000000000c8973d);
sram_add_entry(0, 1, 2132, 4, 128'h40200000000000000000063403b);
sram_add_entry(0, 1, 2136, 4, 128'h4020000000000000000003b10ba);
sram_add_entry(0, 1, 2140, 4, 128'h4020000000000000000002ce7ba);
sram_add_entry(0, 1, 2144, 4, 128'h40200000000000000000000ea87);
sram_add_entry(0, 1, 2148, 4, 128'h40200000000000000000050badf);
sram_add_entry(0, 1, 2152, 4, 128'h4020000000000000000005b2fbb);
sram_add_entry(0, 1, 2156, 4, 128'h402000000000000000000ac32d9);
sram_add_entry(0, 1, 2160, 4, 128'h402000000000000000000175207);
sram_add_entry(0, 1, 2164, 4, 128'h402000000000000000000ce27f9);
sram_add_entry(0, 1, 2168, 4, 128'h40200000000000000000075d740);
sram_add_entry(0, 1, 2172, 4, 128'h40200000000000000000076d79a);
sram_add_entry(0, 1, 2176, 4, 128'h4020000000000000000007390f8);
sram_add_entry(0, 1, 2180, 4, 128'h402000000000000000000b963bf);
sram_add_entry(0, 1, 2184, 4, 128'h402000000000000000000026405);
sram_add_entry(0, 1, 2188, 4, 128'h402000000000000000000a04b21);
sram_add_entry(0, 1, 2192, 4, 128'h402000000000000000000a30541);
sram_add_entry(0, 1, 2196, 4, 128'h4020000000000000000008927b6);
sram_add_entry(0, 1, 2200, 4, 128'h4020000000000000000009cc1c0);
sram_add_entry(0, 1, 2204, 4, 128'h4020000000000000000003ba3f5);
sram_add_entry(0, 1, 2208, 4, 128'h402000000000000000000352e1d);
sram_add_entry(0, 1, 2212, 4, 128'h402000000000000000000c2fbc1);
sram_add_entry(0, 1, 2216, 4, 128'h4020000000000000000004cbb09);
sram_add_entry(0, 1, 2220, 4, 128'h402000000000000000000ffbbbf);
sram_add_entry(0, 1, 2224, 4, 128'h402000000000000000000b682c8);
sram_add_entry(0, 1, 2228, 4, 128'h40200000000000000000052c4da);
sram_add_entry(0, 1, 2232, 4, 128'h402000000000000000000312a41);
sram_add_entry(0, 1, 2236, 4, 128'h40200000000000000000008b4d5);
sram_add_entry(0, 1, 2240, 4, 128'h402000000000000000000f3a2ad);
sram_add_entry(0, 1, 2244, 4, 128'h4020000000000000000006e7c4f);
sram_add_entry(0, 1, 2248, 4, 128'h402000000000000000000ded8dc);
sram_add_entry(0, 1, 2252, 4, 128'h40200000000000000000001dc81);
sram_add_entry(0, 1, 2256, 4, 128'h4020000000000000000000fbaf9);
sram_add_entry(0, 1, 2260, 4, 128'h40200000000000000000061584b);
sram_add_entry(0, 1, 2264, 4, 128'h4020000000000000000007649b8);
sram_add_entry(0, 1, 2268, 4, 128'h4020000000000000000005f5cd1);
sram_add_entry(0, 1, 2272, 4, 128'h402000000000000000000f10131);
sram_add_entry(0, 1, 2276, 4, 128'h40200000000000000000072671c);
sram_add_entry(0, 1, 2280, 4, 128'h402000000000000000000d3785d);
sram_add_entry(0, 1, 2284, 4, 128'h402000000000000000000a29593);
sram_add_entry(0, 1, 2288, 4, 128'h402000000000000000000954c60);
sram_add_entry(0, 1, 2292, 4, 128'h402000000000000000000c17e8e);
sram_add_entry(0, 1, 2296, 4, 128'h40200000000000000000009a7ba);
sram_add_entry(0, 1, 2300, 4, 128'h4020000000000000000007072f3);
sram_add_entry(0, 1, 2304, 4, 128'h40200000000000000000078fcbf);
sram_add_entry(0, 1, 2308, 4, 128'h40200000000000000000043c1b7);
sram_add_entry(0, 1, 2312, 4, 128'h402000000000000000000b08007);
sram_add_entry(0, 1, 2316, 4, 128'h402000000000000000000150566);
sram_add_entry(0, 1, 2320, 4, 128'h402000000000000000000a9a978);
sram_add_entry(0, 1, 2324, 4, 128'h402000000000000000000c86b86);
sram_add_entry(0, 1, 2328, 4, 128'h402000000000000000000f6a9b4);
sram_add_entry(0, 1, 2332, 4, 128'h402000000000000000000bd5e1d);
sram_add_entry(0, 1, 2336, 4, 128'h4020000000000000000006bdf3d);
sram_add_entry(0, 1, 2340, 4, 128'h4020000000000000000008848ec);
sram_add_entry(0, 1, 2344, 4, 128'h4020000000000000000002de4cb);
sram_add_entry(0, 1, 2348, 4, 128'h402000000000000000000729081);
sram_add_entry(0, 1, 2352, 4, 128'h4020000000000000000006a8d3d);
sram_add_entry(0, 1, 2356, 4, 128'h402000000000000000000b986e7);
sram_add_entry(0, 1, 2360, 4, 128'h40200000000000000000053a9dc);
sram_add_entry(0, 1, 2364, 4, 128'h402000000000000000000495aab);
sram_add_entry(0, 1, 2368, 4, 128'h4020000000000000000002243c5);
sram_add_entry(0, 1, 2372, 4, 128'h402000000000000000000932bc5);
sram_add_entry(0, 1, 2376, 4, 128'h402000000000000000000c7e5a1);
sram_add_entry(0, 1, 2380, 4, 128'h402000000000000000000519f51);
sram_add_entry(0, 1, 2384, 4, 128'h40200000000000000000031d9d3);
sram_add_entry(0, 1, 2388, 4, 128'h4020000000000000000006c648c);
sram_add_entry(0, 1, 2392, 4, 128'h402000000000000000000ca4098);
sram_add_entry(0, 1, 2396, 4, 128'h402000000000000000000e6aa63);
sram_add_entry(0, 1, 2400, 4, 128'h4020000000000000000009898d6);
sram_add_entry(0, 1, 2404, 4, 128'h4020000000000000000002e0ee6);
sram_add_entry(0, 1, 2408, 4, 128'h4020000000000000000007de959);
sram_add_entry(0, 1, 2412, 4, 128'h40200000000000000000022ed5e);
sram_add_entry(0, 1, 2416, 4, 128'h402000000000000000000ef9cd4);
sram_add_entry(0, 1, 2420, 4, 128'h4020000000000000000009e573b);
sram_add_entry(0, 1, 2424, 4, 128'h402000000000000000000a4a6bf);
sram_add_entry(0, 1, 2428, 4, 128'h40200000000000000000096fae7);
sram_add_entry(0, 1, 2432, 4, 128'h402000000000000000000cdbaec);
sram_add_entry(0, 1, 2436, 4, 128'h402000000000000000000f9a463);
sram_add_entry(0, 1, 2440, 4, 128'h4020000000000000000004e36e0);
sram_add_entry(0, 1, 2444, 4, 128'h402000000000000000000f0a7a9);
sram_add_entry(0, 1, 2448, 4, 128'h4020000000000000000001ae7e7);
sram_add_entry(0, 1, 2452, 4, 128'h402000000000000000000facdcc);
sram_add_entry(0, 1, 2456, 4, 128'h402000000000000000000057f90);
sram_add_entry(0, 1, 2460, 4, 128'h402000000000000000000b782da);
sram_add_entry(0, 1, 2464, 4, 128'h4020000000000000000000068b3);
sram_add_entry(0, 1, 2468, 4, 128'h4020000000000000000003a8542);
sram_add_entry(0, 1, 2472, 4, 128'h402000000000000000000662a36);
sram_add_entry(0, 1, 2476, 4, 128'h402000000000000000000c447e7);
sram_add_entry(0, 1, 2480, 4, 128'h402000000000000000000428275);
sram_add_entry(0, 1, 2484, 4, 128'h402000000000000000000207e9f);
sram_add_entry(0, 1, 2488, 4, 128'h402000000000000000000b5de9b);
sram_add_entry(0, 1, 2492, 4, 128'h402000000000000000000bdfb18);
sram_add_entry(0, 1, 2496, 4, 128'h4020000000000000000003a7a85);
sram_add_entry(0, 1, 2500, 4, 128'h4020000000000000000006b085d);
sram_add_entry(0, 1, 2504, 4, 128'h402000000000000000000e56816);
sram_add_entry(0, 1, 2508, 4, 128'h40200000000000000000018d22b);
sram_add_entry(0, 1, 2512, 4, 128'h402000000000000000000fd73c1);
sram_add_entry(0, 1, 2516, 4, 128'h402000000000000000000f65166);
sram_add_entry(0, 1, 2520, 4, 128'h402000000000000000000aea4f6);
sram_add_entry(0, 1, 2524, 4, 128'h402000000000000000000378ad7);
sram_add_entry(0, 1, 2528, 4, 128'h4020000000000000000007215cb);
sram_add_entry(0, 1, 2532, 4, 128'h4020000000000000000004370d3);
sram_add_entry(0, 1, 2536, 4, 128'h402000000000000000000e0bb48);
sram_add_entry(0, 1, 2540, 4, 128'h402000000000000000000dd2dbc);
sram_add_entry(0, 1, 2544, 4, 128'h402000000000000000000d10c0d);
sram_add_entry(0, 1, 2548, 4, 128'h40200000000000000000045ca7b);
sram_add_entry(0, 1, 2552, 4, 128'h40200000000000000000050ec64);
sram_add_entry(0, 1, 2556, 4, 128'h402000000000000000000906144);
sram_add_entry(0, 1, 2560, 4, 128'h402000000000000000000112dc1);
sram_add_entry(0, 1, 2564, 4, 128'h4020000000000000000005b36ae);
sram_add_entry(0, 1, 2568, 4, 128'h4020000000000000000006a5c37);
sram_add_entry(0, 1, 2572, 4, 128'h40200000000000000000024a942);
sram_add_entry(0, 1, 2576, 4, 128'h402000000000000000000048e2b);
sram_add_entry(0, 1, 2580, 4, 128'h40200000000000000000077fa27);
sram_add_entry(0, 1, 2584, 4, 128'h40200000000000000000078b151);
sram_add_entry(0, 1, 2588, 4, 128'h402000000000000000000a47604);
sram_add_entry(0, 1, 2592, 4, 128'h402000000000000000000594a3f);
sram_add_entry(0, 1, 2596, 4, 128'h402000000000000000000af2e91);
sram_add_entry(0, 1, 2600, 4, 128'h40200000000000000000054f406);
sram_add_entry(0, 1, 2604, 4, 128'h402000000000000000000dbd353);
sram_add_entry(0, 1, 2608, 4, 128'h402000000000000000000a961f7);
sram_add_entry(0, 1, 2612, 4, 128'h402000000000000000000655384);
sram_add_entry(0, 1, 2616, 4, 128'h40200000000000000000001b8b2);
sram_add_entry(0, 1, 2620, 4, 128'h402000000000000000000b646a0);
sram_add_entry(0, 1, 2624, 4, 128'h402000000000000000000c35541);
sram_add_entry(0, 1, 2628, 4, 128'h402000000000000000000aa459d);
sram_add_entry(0, 1, 2632, 4, 128'h402000000000000000000759b4f);
sram_add_entry(0, 1, 2636, 4, 128'h40200000000000000000010b764);
sram_add_entry(0, 1, 2640, 4, 128'h4020000000000000000007f2ca2);
sram_add_entry(0, 1, 2644, 4, 128'h402000000000000000000009605);
sram_add_entry(0, 1, 2648, 4, 128'h402000000000000000000880ee7);
sram_add_entry(0, 1, 2652, 4, 128'h402000000000000000000eced99);
sram_add_entry(0, 1, 2656, 4, 128'h4020000000000000000008a05ca);
sram_add_entry(0, 1, 2660, 4, 128'h40200000000000000000066baf9);
sram_add_entry(0, 1, 2664, 4, 128'h40200000000000000000096805d);
sram_add_entry(0, 1, 2668, 4, 128'h4020000000000000000000e3de2);
sram_add_entry(0, 1, 2672, 4, 128'h40200000000000000000015e3df);
sram_add_entry(0, 1, 2676, 4, 128'h402000000000000000000a47712);
sram_add_entry(0, 1, 2680, 4, 128'h4020000000000000000001932f3);
sram_add_entry(0, 1, 2684, 4, 128'h40200000000000000000015d54c);
sram_add_entry(0, 1, 2688, 4, 128'h4020000000000000000008e6097);
sram_add_entry(0, 1, 2692, 4, 128'h402000000000000000000026723);
sram_add_entry(0, 1, 2696, 4, 128'h4020000000000000000002d4201);
sram_add_entry(0, 1, 2700, 4, 128'h40200000000000000000064a019);
sram_add_entry(0, 1, 2704, 4, 128'h402000000000000000000052068);
sram_add_entry(0, 1, 2708, 4, 128'h4020000000000000000004fc87f);
sram_add_entry(0, 1, 2712, 4, 128'h402000000000000000000354c4a);
sram_add_entry(0, 1, 2716, 4, 128'h402000000000000000000c084df);
sram_add_entry(0, 1, 2720, 4, 128'h402000000000000000000e3af6c);
sram_add_entry(0, 1, 2724, 4, 128'h4020000000000000000009b4c6a);
sram_add_entry(0, 1, 2728, 4, 128'h4020000000000000000004fe061);
sram_add_entry(0, 1, 2732, 4, 128'h402000000000000000000668b54);
sram_add_entry(0, 1, 2736, 4, 128'h402000000000000000000b7d2fa);
sram_add_entry(0, 1, 2740, 4, 128'h4020000000000000000007b394b);
sram_add_entry(0, 1, 2744, 4, 128'h402000000000000000000a0d693);
sram_add_entry(0, 1, 2748, 4, 128'h402000000000000000000ecb9e8);
sram_add_entry(0, 1, 2752, 4, 128'h402000000000000000000fa6dcb);
sram_add_entry(0, 1, 2756, 4, 128'h402000000000000000000549727);
sram_add_entry(0, 1, 2760, 4, 128'h402000000000000000000563be7);
sram_add_entry(0, 1, 2764, 4, 128'h402000000000000000000efc0f2);
sram_add_entry(0, 1, 2768, 4, 128'h402000000000000000000c5e4f2);
sram_add_entry(0, 1, 2772, 4, 128'h40200000000000000000097e2e2);
sram_add_entry(0, 1, 2776, 4, 128'h402000000000000000000d71d42);
sram_add_entry(0, 1, 2780, 4, 128'h4020000000000000000002cc08f);
sram_add_entry(0, 1, 2784, 4, 128'h4020000000000000000006e18f9);
sram_add_entry(0, 1, 2788, 4, 128'h4020000000000000000000fdf59);
sram_add_entry(0, 1, 2792, 4, 128'h4020000000000000000008f22b0);
sram_add_entry(0, 1, 2796, 4, 128'h402000000000000000000f70e50);
sram_add_entry(0, 1, 2800, 4, 128'h40200000000000000000065c364);
sram_add_entry(0, 0, 0, 4, 128'h7ab000000000000000000deadbf);
sram_add_entry(0, 0, 4, 4, 128'h4020000000000000000007f1ea9);
sram_add_entry(0, 0, 8, 4, 128'h40200000000000000000018d7d4);
sram_add_entry(0, 0, 12, 4, 128'h402000000000000000000879503);
sram_add_entry(0, 0, 16, 4, 128'h402000000000000000000795e9d);
sram_add_entry(0, 0, 20, 4, 128'h402000000000000000000d8811f);
sram_add_entry(0, 0, 24, 4, 128'h402000000000000000000f72c4f);
sram_add_entry(0, 0, 28, 4, 128'h40200000000000000000045bc37);
sram_add_entry(0, 0, 32, 4, 128'h402000000000000000000a9ca1e);
sram_add_entry(0, 0, 36, 4, 128'h40200000000000000000095fadc);
sram_add_entry(0, 0, 40, 4, 128'h402000000000000000000fd7856);
sram_add_entry(0, 0, 44, 4, 128'h4020000000000000000003ac1d0);
sram_add_entry(0, 0, 48, 4, 128'h4020000000000000000000c47e0);
sram_add_entry(0, 0, 52, 4, 128'h402000000000000000000fb27f9);
sram_add_entry(0, 0, 56, 4, 128'h40200000000000000000018fca4);
sram_add_entry(0, 0, 60, 4, 128'h4020000000000000000002e4356);
sram_add_entry(0, 0, 64, 4, 128'h40200000000000000000056a40c);
sram_add_entry(0, 0, 68, 4, 128'h40200000000000000000018540e);
sram_add_entry(0, 0, 72, 4, 128'h402000000000000000000ea2b44);
sram_add_entry(0, 0, 76, 4, 128'h40200000000000000000084c769);
sram_add_entry(0, 0, 80, 4, 128'h4020000000000000000009ae0b9);
sram_add_entry(0, 0, 84, 4, 128'h402000000000000000000a15356);
sram_add_entry(0, 0, 88, 4, 128'h4020000000000000000005a0605);
sram_add_entry(0, 0, 92, 4, 128'h4020000000000000000006fe0cb);
sram_add_entry(0, 0, 96, 4, 128'h402000000000000000000e646d6);
sram_add_entry(0, 0, 100, 4, 128'h4020000000000000000000a2d6b);
sram_add_entry(0, 0, 104, 4, 128'h402000000000000000000f04d5b);
sram_add_entry(0, 0, 108, 4, 128'h4020000000000000000004c578c);
sram_add_entry(0, 0, 112, 4, 128'h402000000000000000000888d1f);
sram_add_entry(0, 0, 116, 4, 128'h4020000000000000000002ca3fe);
sram_add_entry(0, 0, 120, 4, 128'h40200000000000000000063455b);
sram_add_entry(0, 0, 124, 4, 128'h4020000000000000000002768c3);
sram_add_entry(0, 0, 128, 4, 128'h4020000000000000000007cb8cb);
sram_add_entry(0, 0, 132, 4, 128'h40200000000000000000062f735);
sram_add_entry(0, 0, 136, 4, 128'h4020000000000000000002fa2ac);
sram_add_entry(0, 0, 140, 4, 128'h4020000000000000000006b0b30);
sram_add_entry(0, 0, 144, 4, 128'h402000000000000000000dc4120);
sram_add_entry(0, 0, 148, 4, 128'h402000000000000000000d471aa);
sram_add_entry(0, 0, 152, 4, 128'h40200000000000000000040a7fc);
sram_add_entry(0, 0, 156, 4, 128'h402000000000000000000ac33c6);
sram_add_entry(0, 0, 160, 4, 128'h402000000000000000000109775);
sram_add_entry(0, 0, 164, 4, 128'h402000000000000000000c3ff40);
sram_add_entry(0, 0, 168, 4, 128'h402000000000000000000283e24);
sram_add_entry(0, 0, 172, 4, 128'h402000000000000000000d2bca2);
sram_add_entry(0, 0, 176, 4, 128'h4020000000000000000005178a5);
sram_add_entry(0, 0, 180, 4, 128'h4020000000000000000009ab1a5);
sram_add_entry(0, 0, 184, 4, 128'h402000000000000000000dd0418);
sram_add_entry(0, 0, 188, 4, 128'h4020000000000000000004341e8);
sram_add_entry(0, 0, 192, 4, 128'h402000000000000000000beafd2);
sram_add_entry(0, 0, 196, 4, 128'h402000000000000000000653c68);
sram_add_entry(0, 0, 200, 4, 128'h402000000000000000000c2f7fb);
sram_add_entry(0, 0, 204, 4, 128'h4020000000000000000002ec425);
sram_add_entry(0, 0, 208, 4, 128'h40200000000000000000039f1b8);
sram_add_entry(0, 0, 212, 4, 128'h40200000000000000000065b81f);
sram_add_entry(0, 0, 216, 4, 128'h402000000000000000000e84bff);
sram_add_entry(0, 0, 220, 4, 128'h4020000000000000000006f12c1);
sram_add_entry(0, 0, 224, 4, 128'h402000000000000000000638539);
sram_add_entry(0, 0, 228, 4, 128'h40200000000000000000074386b);
sram_add_entry(0, 0, 232, 4, 128'h4020000000000000000006ec296);
sram_add_entry(0, 0, 236, 4, 128'h4020000000000000000009dc45a);
sram_add_entry(0, 0, 240, 4, 128'h4020000000000000000007bdeb2);
sram_add_entry(0, 0, 244, 4, 128'h402000000000000000000109400);
sram_add_entry(0, 0, 248, 4, 128'h4020000000000000000003ed34b);
sram_add_entry(0, 0, 252, 4, 128'h40200000000000000000083a39a);
sram_add_entry(0, 0, 256, 4, 128'h402000000000000000000b39350);
sram_add_entry(0, 0, 260, 4, 128'h4020000000000000000003fd68e);
sram_add_entry(0, 0, 264, 4, 128'h402000000000000000000168dc8);
sram_add_entry(0, 0, 268, 4, 128'h402000000000000000000c7d864);
sram_add_entry(0, 0, 272, 4, 128'h4020000000000000000006ac4b8);
sram_add_entry(0, 0, 276, 4, 128'h40200000000000000000029c5fa);
sram_add_entry(0, 0, 280, 4, 128'h4020000000000000000007775e4);
sram_add_entry(0, 0, 284, 4, 128'h402000000000000000000354a38);
sram_add_entry(0, 0, 288, 4, 128'h402000000000000000000482f82);
sram_add_entry(0, 0, 292, 4, 128'h4020000000000000000008f4dc7);
sram_add_entry(0, 0, 296, 4, 128'h4020000000000000000002f794e);
sram_add_entry(0, 0, 300, 4, 128'h402000000000000000000c688bd);
sram_add_entry(0, 0, 304, 4, 128'h4020000000000000000008c6bf8);
sram_add_entry(0, 0, 308, 4, 128'h4020000000000000000004a580d);
sram_add_entry(0, 0, 312, 4, 128'h402000000000000000000e51d07);
sram_add_entry(0, 0, 316, 4, 128'h4020000000000000000006576cb);
sram_add_entry(0, 0, 320, 4, 128'h402000000000000000000672b33);
sram_add_entry(0, 0, 324, 4, 128'h402000000000000000000765369);
sram_add_entry(0, 0, 328, 4, 128'h402000000000000000000065548);
sram_add_entry(0, 0, 332, 4, 128'h402000000000000000000fa8b7f);
sram_add_entry(0, 0, 336, 4, 128'h4020000000000000000009e0149);
sram_add_entry(0, 0, 340, 4, 128'h4020000000000000000003700bc);
sram_add_entry(0, 0, 344, 4, 128'h402000000000000000000a26d54);
sram_add_entry(0, 0, 348, 4, 128'h402000000000000000000485e50);
sram_add_entry(0, 0, 352, 4, 128'h4020000000000000000004e377c);
sram_add_entry(0, 0, 356, 4, 128'h402000000000000000000290bd8);
sram_add_entry(0, 0, 360, 4, 128'h40200000000000000000079eac3);
sram_add_entry(0, 0, 364, 4, 128'h402000000000000000000aeb963);
sram_add_entry(0, 0, 368, 4, 128'h4020000000000000000000e60f6);
sram_add_entry(0, 0, 372, 4, 128'h402000000000000000000ebc64c);
sram_add_entry(0, 0, 376, 4, 128'h402000000000000000000fd79da);
sram_add_entry(0, 0, 380, 4, 128'h4020000000000000000005f903f);
sram_add_entry(0, 0, 384, 4, 128'h4020000000000000000008c6098);
sram_add_entry(0, 0, 388, 4, 128'h40200000000000000000052bbf8);
sram_add_entry(0, 0, 392, 4, 128'h40200000000000000000067064a);
sram_add_entry(0, 0, 396, 4, 128'h402000000000000000000eda0ac);
sram_add_entry(0, 0, 400, 4, 128'h4020000000000000000009fe0b2);
sram_add_entry(0, 0, 404, 4, 128'h4020000000000000000002b0b9e);
sram_add_entry(0, 0, 408, 4, 128'h4020000000000000000008ed315);
sram_add_entry(0, 0, 412, 4, 128'h4020000000000000000003fa5eb);
sram_add_entry(0, 0, 416, 4, 128'h402000000000000000000d5a9ea);
sram_add_entry(0, 0, 420, 4, 128'h4020000000000000000003b5063);
sram_add_entry(0, 0, 424, 4, 128'h4020000000000000000003de498);
sram_add_entry(0, 0, 428, 4, 128'h40200000000000000000034d05b);
sram_add_entry(0, 0, 432, 4, 128'h4020000000000000000009906b4);
sram_add_entry(0, 0, 436, 4, 128'h4020000000000000000008e8559);
sram_add_entry(0, 0, 440, 4, 128'h4020000000000000000000e3f52);
sram_add_entry(0, 0, 444, 4, 128'h4020000000000000000004b4571);
sram_add_entry(0, 0, 448, 4, 128'h4020000000000000000001da95e);
sram_add_entry(0, 0, 452, 4, 128'h402000000000000000000f8a77d);
sram_add_entry(0, 0, 456, 4, 128'h4020000000000000000000773e7);
sram_add_entry(0, 0, 460, 4, 128'h402000000000000000000cc18d8);
sram_add_entry(0, 0, 464, 4, 128'h402000000000000000000523f2c);
sram_add_entry(0, 0, 468, 4, 128'h402000000000000000000d32eb1);
sram_add_entry(0, 0, 472, 4, 128'h402000000000000000000b10a04);
sram_add_entry(0, 0, 476, 4, 128'h4020000000000000000009e289a);
sram_add_entry(0, 0, 480, 4, 128'h4020000000000000000003f745c);
sram_add_entry(0, 0, 484, 4, 128'h402000000000000000000b4d716);
sram_add_entry(0, 0, 488, 4, 128'h402000000000000000000353aba);
sram_add_entry(0, 0, 492, 4, 128'h402000000000000000000138266);
sram_add_entry(0, 0, 496, 4, 128'h40200000000000000000098c3a8);
sram_add_entry(0, 0, 500, 4, 128'h402000000000000000000a72bb0);
sram_add_entry(0, 0, 504, 4, 128'h402000000000000000000f0a808);
sram_add_entry(0, 0, 508, 4, 128'h4020000000000000000002ecc7c);
sram_add_entry(0, 0, 512, 4, 128'h40200000000000000000070432e);
sram_add_entry(0, 0, 516, 4, 128'h4020000000000000000009e5629);
sram_add_entry(0, 0, 520, 4, 128'h402000000000000000000b9028f);
sram_add_entry(0, 0, 524, 4, 128'h4020000000000000000007d192f);
sram_add_entry(0, 0, 528, 4, 128'h4020000000000000000009f9291);
sram_add_entry(0, 0, 532, 4, 128'h402000000000000000000ee6a20);
sram_add_entry(0, 0, 536, 4, 128'h40200000000000000000053672d);
sram_add_entry(0, 0, 540, 4, 128'h402000000000000000000dd027c);
sram_add_entry(0, 0, 544, 4, 128'h4020000000000000000000dc08c);
sram_add_entry(0, 0, 548, 4, 128'h40200000000000000000058402c);
sram_add_entry(0, 0, 552, 4, 128'h402000000000000000000c81a4a);
sram_add_entry(0, 0, 556, 4, 128'h402000000000000000000edd5d3);
sram_add_entry(0, 0, 560, 4, 128'h402000000000000000000004b52);
sram_add_entry(0, 0, 564, 4, 128'h402000000000000000000e03ed4);
sram_add_entry(0, 0, 568, 4, 128'h4020000000000000000007e9436);
sram_add_entry(0, 0, 572, 4, 128'h402000000000000000000784bef);
sram_add_entry(0, 0, 576, 4, 128'h40200000000000000000042f39d);
sram_add_entry(0, 0, 580, 4, 128'h402000000000000000000be6a7e);
sram_add_entry(0, 0, 584, 4, 128'h402000000000000000000826f57);
sram_add_entry(0, 0, 588, 4, 128'h402000000000000000000029e2c);
sram_add_entry(0, 0, 592, 4, 128'h40200000000000000000029c960);
sram_add_entry(0, 0, 596, 4, 128'h40200000000000000000019c756);
sram_add_entry(0, 0, 600, 4, 128'h40200000000000000000001fbdf);
sram_add_entry(0, 0, 604, 4, 128'h4020000000000000000000798a3);
sram_add_entry(0, 0, 608, 4, 128'h402000000000000000000376c99);
sram_add_entry(0, 0, 612, 4, 128'h4020000000000000000002e7c93);
sram_add_entry(0, 0, 616, 4, 128'h4020000000000000000006e0c48);
sram_add_entry(0, 0, 620, 4, 128'h4020000000000000000007848e4);
sram_add_entry(0, 0, 624, 4, 128'h402000000000000000000eab49b);
sram_add_entry(0, 0, 628, 4, 128'h4020000000000000000003c4183);
sram_add_entry(0, 0, 632, 4, 128'h402000000000000000000206e77);
sram_add_entry(0, 0, 636, 4, 128'h40200000000000000000060af7b);
sram_add_entry(0, 0, 640, 4, 128'h402000000000000000000532847);
sram_add_entry(0, 0, 644, 4, 128'h402000000000000000000bad608);
sram_add_entry(0, 0, 648, 4, 128'h40200000000000000000047a19a);
sram_add_entry(0, 0, 652, 4, 128'h402000000000000000000f8c422);
sram_add_entry(0, 0, 656, 4, 128'h4020000000000000000009c50ab);
sram_add_entry(0, 0, 660, 4, 128'h4020000000000000000002c4a16);
sram_add_entry(0, 0, 664, 4, 128'h402000000000000000000e2f212);
sram_add_entry(0, 0, 668, 4, 128'h40200000000000000000032b6e2);
sram_add_entry(0, 0, 672, 4, 128'h402000000000000000000501cd9);
sram_add_entry(0, 0, 676, 4, 128'h40200000000000000000059d817);
sram_add_entry(0, 0, 680, 4, 128'h40200000000000000000079c4b3);
sram_add_entry(0, 0, 684, 4, 128'h402000000000000000000dbfb38);
sram_add_entry(0, 0, 688, 4, 128'h4020000000000000000003c8d91);
sram_add_entry(0, 0, 692, 4, 128'h402000000000000000000700b97);
sram_add_entry(0, 0, 696, 4, 128'h4020000000000000000006a6798);
sram_add_entry(0, 0, 700, 4, 128'h402000000000000000000b16541);
sram_add_entry(0, 0, 704, 4, 128'h402000000000000000000148fdc);
sram_add_entry(0, 0, 708, 4, 128'h402000000000000000000c77ae0);
sram_add_entry(0, 0, 712, 4, 128'h402000000000000000000289a41);
sram_add_entry(0, 0, 716, 4, 128'h402000000000000000000cce9c6);
sram_add_entry(0, 0, 720, 4, 128'h4020000000000000000003293d0);
sram_add_entry(0, 0, 724, 4, 128'h40200000000000000000085fe27);
sram_add_entry(0, 0, 728, 4, 128'h4020000000000000000007de321);
sram_add_entry(0, 0, 732, 4, 128'h402000000000000000000556878);
sram_add_entry(0, 0, 736, 4, 128'h402000000000000000000a2e200);
sram_add_entry(0, 0, 740, 4, 128'h402000000000000000000f7b199);
sram_add_entry(0, 0, 744, 4, 128'h4020000000000000000004e7d0f);
sram_add_entry(0, 0, 748, 4, 128'h4020000000000000000002932d5);
sram_add_entry(0, 0, 752, 4, 128'h402000000000000000000f10ee2);
sram_add_entry(0, 0, 756, 4, 128'h402000000000000000000d3cb30);
sram_add_entry(0, 0, 760, 4, 128'h402000000000000000000dc4082);
sram_add_entry(0, 0, 764, 4, 128'h4020000000000000000004680df);
sram_add_entry(0, 0, 768, 4, 128'h4020000000000000000003e3ace);
sram_add_entry(0, 0, 772, 4, 128'h402000000000000000000278237);
sram_add_entry(0, 0, 776, 4, 128'h402000000000000000000f58b4b);
sram_add_entry(0, 0, 780, 4, 128'h40200000000000000000053a60b);
sram_add_entry(0, 0, 784, 4, 128'h40200000000000000000029bce4);
sram_add_entry(0, 0, 788, 4, 128'h402000000000000000000bf1a0a);
sram_add_entry(0, 0, 792, 4, 128'h402000000000000000000e19318);
sram_add_entry(0, 0, 796, 4, 128'h40200000000000000000044d266);
sram_add_entry(0, 0, 800, 4, 128'h402000000000000000000a6b455);
sram_add_entry(0, 0, 804, 4, 128'h402000000000000000000a1ed9d);
sram_add_entry(0, 0, 808, 4, 128'h4020000000000000000004fc0f7);
sram_add_entry(0, 0, 812, 4, 128'h40200000000000000000083eaaf);
sram_add_entry(0, 0, 816, 4, 128'h40200000000000000000001d8f2);
sram_add_entry(0, 0, 820, 4, 128'h4020000000000000000000c8461);
sram_add_entry(0, 0, 824, 4, 128'h4020000000000000000005a9ad8);
sram_add_entry(0, 0, 828, 4, 128'h40200000000000000000045adc4);
sram_add_entry(0, 0, 832, 4, 128'h40200000000000000000044e7f5);
sram_add_entry(0, 0, 836, 4, 128'h4020000000000000000004a5dba);
sram_add_entry(0, 0, 840, 4, 128'h40200000000000000000082d37a);
sram_add_entry(0, 0, 844, 4, 128'h402000000000000000000a5936e);
sram_add_entry(0, 0, 848, 4, 128'h40200000000000000000007b239);
sram_add_entry(0, 0, 852, 4, 128'h40200000000000000000012fd45);
sram_add_entry(0, 0, 856, 4, 128'h402000000000000000000842ec1);
sram_add_entry(0, 0, 860, 4, 128'h4020000000000000000005fee07);
sram_add_entry(0, 0, 864, 4, 128'h402000000000000000000386dc0);
sram_add_entry(0, 0, 868, 4, 128'h40200000000000000000030a003);
sram_add_entry(0, 0, 872, 4, 128'h40200000000000000000069dabf);
sram_add_entry(0, 0, 876, 4, 128'h4020000000000000000000c8cd9);
sram_add_entry(0, 0, 880, 4, 128'h40200000000000000000020926d);
sram_add_entry(0, 0, 884, 4, 128'h402000000000000000000c358af);
sram_add_entry(0, 0, 888, 4, 128'h4020000000000000000005bb9eb);
sram_add_entry(0, 0, 892, 4, 128'h402000000000000000000b1e73e);
sram_add_entry(0, 0, 896, 4, 128'h402000000000000000000591f46);
sram_add_entry(0, 0, 900, 4, 128'h4020000000000000000007367d3);
sram_add_entry(0, 0, 904, 4, 128'h402000000000000000000638b62);
sram_add_entry(0, 0, 908, 4, 128'h402000000000000000000637b90);
sram_add_entry(0, 0, 912, 4, 128'h4020000000000000000008d74b6);
sram_add_entry(0, 0, 916, 4, 128'h4020000000000000000005c8f52);
sram_add_entry(0, 0, 920, 4, 128'h402000000000000000000d7ee49);
sram_add_entry(0, 0, 924, 4, 128'h402000000000000000000d72b91);
sram_add_entry(0, 0, 928, 4, 128'h402000000000000000000816c24);
sram_add_entry(0, 0, 932, 4, 128'h402000000000000000000de97a8);
sram_add_entry(0, 0, 936, 4, 128'h4020000000000000000004ef26b);
sram_add_entry(0, 0, 940, 4, 128'h402000000000000000000afbc7c);
sram_add_entry(0, 0, 944, 4, 128'h402000000000000000000337d7d);
sram_add_entry(0, 0, 948, 4, 128'h402000000000000000000781a2b);
sram_add_entry(0, 0, 952, 4, 128'h402000000000000000000b4e99c);
sram_add_entry(0, 0, 956, 4, 128'h402000000000000000000a1d931);
sram_add_entry(0, 0, 960, 4, 128'h4020000000000000000002e3027);
sram_add_entry(0, 0, 964, 4, 128'h402000000000000000000f983f9);
sram_add_entry(0, 0, 968, 4, 128'h40200000000000000000056ed80);
sram_add_entry(0, 0, 972, 4, 128'h4020000000000000000005200ab);
sram_add_entry(0, 0, 976, 4, 128'h402000000000000000000637797);
sram_add_entry(0, 0, 980, 4, 128'h402000000000000000000dd2137);
sram_add_entry(0, 0, 984, 4, 128'h402000000000000000000fd2416);
sram_add_entry(0, 0, 988, 4, 128'h402000000000000000000f3a4f0);
sram_add_entry(0, 0, 992, 4, 128'h40200000000000000000044c886);
sram_add_entry(0, 0, 996, 4, 128'h402000000000000000000ceb410);
sram_add_entry(0, 0, 1000, 4, 128'h402000000000000000000f59b12);
sram_add_entry(0, 0, 1004, 4, 128'h402000000000000000000e49bd0);
sram_add_entry(0, 0, 1008, 4, 128'h402000000000000000000638997);
sram_add_entry(0, 0, 1012, 4, 128'h4020000000000000000002f7580);
sram_add_entry(0, 0, 1016, 4, 128'h4020000000000000000001c10a8);
sram_add_entry(0, 0, 1020, 4, 128'h402000000000000000000879f04);
sram_add_entry(0, 0, 1024, 4, 128'h402000000000000000000bab2c4);
sram_add_entry(0, 0, 1028, 4, 128'h402000000000000000000a22715);
sram_add_entry(0, 0, 1032, 4, 128'h402000000000000000000f23b5e);
sram_add_entry(0, 0, 1036, 4, 128'h402000000000000000000fdc001);
sram_add_entry(0, 0, 1040, 4, 128'h402000000000000000000288bf0);
sram_add_entry(0, 0, 1044, 4, 128'h402000000000000000000662d40);
sram_add_entry(0, 0, 1048, 4, 128'h40200000000000000000072cef9);
sram_add_entry(0, 0, 1052, 4, 128'h402000000000000000000087666);
sram_add_entry(0, 0, 1056, 4, 128'h402000000000000000000f522c4);
sram_add_entry(0, 0, 1060, 4, 128'h402000000000000000000cf63c5);
sram_add_entry(0, 0, 1064, 4, 128'h402000000000000000000e18e89);
sram_add_entry(0, 0, 1068, 4, 128'h402000000000000000000a2bc46);
sram_add_entry(0, 0, 1072, 4, 128'h40200000000000000000041996f);
sram_add_entry(0, 0, 1076, 4, 128'h4020000000000000000005e2a51);
sram_add_entry(0, 0, 1080, 4, 128'h40200000000000000000046b451);
sram_add_entry(0, 0, 1084, 4, 128'h402000000000000000000ee2aae);
sram_add_entry(0, 0, 1088, 4, 128'h402000000000000000000b33948);
sram_add_entry(0, 0, 1092, 4, 128'h4020000000000000000007587fe);
sram_add_entry(0, 0, 1096, 4, 128'h4020000000000000000004584c5);
sram_add_entry(0, 0, 1100, 4, 128'h4020000000000000000004532c5);
sram_add_entry(0, 0, 1104, 4, 128'h4020000000000000000007754d8);
sram_add_entry(0, 0, 1108, 4, 128'h40200000000000000000002b77b);
sram_add_entry(0, 0, 1112, 4, 128'h4020000000000000000008f7473);
sram_add_entry(0, 0, 1116, 4, 128'h402000000000000000000ff2471);
sram_add_entry(0, 0, 1120, 4, 128'h40200000000000000000014b05f);
sram_add_entry(0, 0, 1124, 4, 128'h402000000000000000000df9570);
sram_add_entry(0, 0, 1128, 4, 128'h402000000000000000000153dbb);
sram_add_entry(0, 0, 1132, 4, 128'h402000000000000000000c5d62c);
sram_add_entry(0, 0, 1136, 4, 128'h4020000000000000000006bf1fb);
sram_add_entry(0, 0, 1140, 4, 128'h40200000000000000000025d7ea);
sram_add_entry(0, 0, 1144, 4, 128'h4020000000000000000007d1082);
sram_add_entry(0, 0, 1148, 4, 128'h4020000000000000000005f39c9);
sram_add_entry(0, 0, 1152, 4, 128'h40200000000000000000009fe99);
sram_add_entry(0, 0, 1156, 4, 128'h4020000000000000000007b04db);
sram_add_entry(0, 0, 1160, 4, 128'h40200000000000000000029dd6a);
sram_add_entry(0, 0, 1164, 4, 128'h4020000000000000000001fcd7e);
sram_add_entry(0, 0, 1168, 4, 128'h4020000000000000000005b635c);
sram_add_entry(0, 0, 1172, 4, 128'h4020000000000000000006eda0f);
sram_add_entry(0, 0, 1176, 4, 128'h402000000000000000000cef008);
sram_add_entry(0, 0, 1180, 4, 128'h40200000000000000000032dc5e);
sram_add_entry(0, 0, 1184, 4, 128'h40200000000000000000050586f);
sram_add_entry(0, 0, 1188, 4, 128'h4020000000000000000006dc367);
sram_add_entry(0, 0, 1192, 4, 128'h4020000000000000000009c1de1);
sram_add_entry(0, 0, 1196, 4, 128'h402000000000000000000fd77d3);
sram_add_entry(0, 0, 1200, 4, 128'h402000000000000000000d3c5d4);
sram_add_entry(0, 0, 1204, 4, 128'h4020000000000000000000fdb0d);
sram_add_entry(0, 0, 1208, 4, 128'h402000000000000000000025d51);
sram_add_entry(0, 0, 1212, 4, 128'h402000000000000000000e88800);
sram_add_entry(0, 0, 1216, 4, 128'h402000000000000000000c08b8e);
sram_add_entry(0, 0, 1220, 4, 128'h4020000000000000000003f0392);
sram_add_entry(0, 0, 1224, 4, 128'h402000000000000000000a02fb5);
sram_add_entry(0, 0, 1228, 4, 128'h40200000000000000000021607f);
sram_add_entry(0, 0, 1232, 4, 128'h4020000000000000000008f612f);
sram_add_entry(0, 0, 1236, 4, 128'h40200000000000000000034a36e);
sram_add_entry(0, 0, 1240, 4, 128'h402000000000000000000899446);
sram_add_entry(0, 0, 1244, 4, 128'h402000000000000000000aeaee1);
sram_add_entry(0, 0, 1248, 4, 128'h4020000000000000000000efa58);
sram_add_entry(0, 0, 1252, 4, 128'h4020000000000000000007c121d);
sram_add_entry(0, 0, 1256, 4, 128'h40200000000000000000084c243);
sram_add_entry(0, 0, 1260, 4, 128'h4020000000000000000006fa6f1);
sram_add_entry(0, 0, 1264, 4, 128'h402000000000000000000e50d93);
sram_add_entry(0, 0, 1268, 4, 128'h40200000000000000000030a2f4);
sram_add_entry(0, 0, 1272, 4, 128'h40200000000000000000028773f);
sram_add_entry(0, 0, 1276, 4, 128'h4020000000000000000000266b7);
sram_add_entry(0, 0, 1280, 4, 128'h402000000000000000000a9817d);
sram_add_entry(0, 0, 1284, 4, 128'h4020000000000000000003920db);
sram_add_entry(0, 0, 1288, 4, 128'h4020000000000000000003bfaad);
sram_add_entry(0, 0, 1292, 4, 128'h402000000000000000000d9c7f1);
sram_add_entry(0, 0, 1296, 4, 128'h4020000000000000000005c0486);
sram_add_entry(0, 0, 1300, 4, 128'h402000000000000000000d00200);
sram_add_entry(0, 0, 1304, 4, 128'h402000000000000000000d49869);
sram_add_entry(0, 0, 1308, 4, 128'h40200000000000000000089ee4e);
sram_add_entry(0, 0, 1312, 4, 128'h402000000000000000000df942f);
sram_add_entry(0, 0, 1316, 4, 128'h40200000000000000000084601d);
sram_add_entry(0, 0, 1320, 4, 128'h4020000000000000000001808be);
sram_add_entry(0, 0, 1324, 4, 128'h402000000000000000000b502fb);
sram_add_entry(0, 0, 1328, 4, 128'h4020000000000000000009f2b20);
sram_add_entry(0, 0, 1332, 4, 128'h402000000000000000000b2fa64);
sram_add_entry(0, 0, 1336, 4, 128'h40200000000000000000080dd3b);
sram_add_entry(0, 0, 1340, 4, 128'h40200000000000000000038568a);
sram_add_entry(0, 0, 1344, 4, 128'h402000000000000000000ea6666);
sram_add_entry(0, 0, 1348, 4, 128'h402000000000000000000dfa001);
sram_add_entry(0, 0, 1352, 4, 128'h4020000000000000000000396ef);
sram_add_entry(0, 0, 1356, 4, 128'h40200000000000000000061ba43);
sram_add_entry(0, 0, 1360, 4, 128'h402000000000000000000080209);
sram_add_entry(0, 0, 1364, 4, 128'h4020000000000000000005b8fa1);
sram_add_entry(0, 0, 1368, 4, 128'h40200000000000000000061c5cc);
sram_add_entry(0, 0, 1372, 4, 128'h402000000000000000000b26ef1);
sram_add_entry(0, 0, 1376, 4, 128'h402000000000000000000407501);
sram_add_entry(0, 0, 1380, 4, 128'h40200000000000000000028ace5);
sram_add_entry(0, 0, 1384, 4, 128'h402000000000000000000c579b9);
sram_add_entry(0, 0, 1388, 4, 128'h4020000000000000000009bfb01);
sram_add_entry(0, 0, 1392, 4, 128'h4020000000000000000000f34eb);
sram_add_entry(0, 0, 1396, 4, 128'h402000000000000000000ab2f3d);
sram_add_entry(0, 0, 1400, 4, 128'h402000000000000000000186408);
sram_add_entry(0, 0, 1404, 4, 128'h40200000000000000000022a3c9);
sram_add_entry(0, 0, 1408, 4, 128'h4020000000000000000009aa041);
sram_add_entry(0, 0, 1412, 4, 128'h402000000000000000000b46f64);
sram_add_entry(0, 0, 1416, 4, 128'h40200000000000000000048548b);
sram_add_entry(0, 0, 1420, 4, 128'h402000000000000000000e7ee30);
sram_add_entry(0, 0, 1424, 4, 128'h4020000000000000000000c7e65);
sram_add_entry(0, 0, 1428, 4, 128'h402000000000000000000c4e05f);
sram_add_entry(0, 0, 1432, 4, 128'h402000000000000000000cdeb94);
sram_add_entry(0, 0, 1436, 4, 128'h402000000000000000000c6fbde);
sram_add_entry(0, 0, 1440, 4, 128'h4020000000000000000004364d2);
sram_add_entry(0, 0, 1444, 4, 128'h40200000000000000000054c878);
sram_add_entry(0, 0, 1448, 4, 128'h402000000000000000000244700);
sram_add_entry(0, 0, 1452, 4, 128'h4020000000000000000003a7f6d);
sram_add_entry(0, 0, 1456, 4, 128'h402000000000000000000e03a58);
sram_add_entry(0, 0, 1460, 4, 128'h402000000000000000000b0efa4);
sram_add_entry(0, 0, 1464, 4, 128'h4020000000000000000001e6831);
sram_add_entry(0, 0, 1468, 4, 128'h402000000000000000000323acf);
sram_add_entry(0, 0, 1472, 4, 128'h4020000000000000000001ab23b);
sram_add_entry(0, 0, 1476, 4, 128'h402000000000000000000153918);
sram_add_entry(0, 0, 1480, 4, 128'h402000000000000000000a376d9);
sram_add_entry(0, 0, 1484, 4, 128'h40200000000000000000066c250);
sram_add_entry(0, 0, 1488, 4, 128'h402000000000000000000f46295);
sram_add_entry(0, 0, 1492, 4, 128'h402000000000000000000909a33);
sram_add_entry(0, 0, 1496, 4, 128'h402000000000000000000b903f6);
sram_add_entry(0, 0, 1500, 4, 128'h402000000000000000000876713);
sram_add_entry(0, 0, 1504, 4, 128'h402000000000000000000f203b1);
sram_add_entry(0, 0, 1508, 4, 128'h4020000000000000000007035e4);
sram_add_entry(0, 0, 1512, 4, 128'h402000000000000000000e24033);
sram_add_entry(0, 0, 1516, 4, 128'h402000000000000000000e8a4a2);
sram_add_entry(0, 0, 1520, 4, 128'h402000000000000000000ece548);
sram_add_entry(0, 0, 1524, 4, 128'h402000000000000000000586dfc);
sram_add_entry(0, 0, 1528, 4, 128'h4020000000000000000008c1319);
sram_add_entry(0, 0, 1532, 4, 128'h402000000000000000000725176);
sram_add_entry(0, 0, 1536, 4, 128'h40200000000000000000056cec2);
sram_add_entry(0, 0, 1540, 4, 128'h402000000000000000000639a04);
sram_add_entry(0, 0, 1544, 4, 128'h4020000000000000000005327e0);
sram_add_entry(0, 0, 1548, 4, 128'h4020000000000000000001462c7);
sram_add_entry(0, 0, 1552, 4, 128'h4020000000000000000000d89f5);
sram_add_entry(0, 0, 1556, 4, 128'h4020000000000000000003902ae);
sram_add_entry(0, 0, 1560, 4, 128'h402000000000000000000a2cbeb);
sram_add_entry(0, 0, 1564, 4, 128'h4020000000000000000000f6681);
sram_add_entry(0, 0, 1568, 4, 128'h4020000000000000000005dcafd);
sram_add_entry(0, 0, 1572, 4, 128'h402000000000000000000691152);
sram_add_entry(0, 0, 1576, 4, 128'h40200000000000000000076bcf7);
sram_add_entry(0, 0, 1580, 4, 128'h402000000000000000000655333);
sram_add_entry(0, 0, 1584, 4, 128'h40200000000000000000067c107);
sram_add_entry(0, 0, 1588, 4, 128'h402000000000000000000bd651c);
sram_add_entry(0, 0, 1592, 4, 128'h402000000000000000000d88fbe);
sram_add_entry(0, 0, 1596, 4, 128'h4020000000000000000003fa26a);
sram_add_entry(0, 0, 1600, 4, 128'h402000000000000000000be3762);
sram_add_entry(0, 0, 1604, 4, 128'h402000000000000000000ee1fc4);
sram_add_entry(0, 0, 1608, 4, 128'h402000000000000000000b30bdf);
sram_add_entry(0, 0, 1612, 4, 128'h402000000000000000000977fec);
sram_add_entry(0, 0, 1616, 4, 128'h402000000000000000000f34eee);
sram_add_entry(0, 0, 1620, 4, 128'h40200000000000000000088c78e);
sram_add_entry(0, 0, 1624, 4, 128'h40200000000000000000050186a);
sram_add_entry(0, 0, 1628, 4, 128'h40200000000000000000022c496);
sram_add_entry(0, 0, 1632, 4, 128'h40200000000000000000074ba14);
sram_add_entry(0, 0, 1636, 4, 128'h4020000000000000000005fa922);
sram_add_entry(0, 0, 1640, 4, 128'h40200000000000000000009f94e);
sram_add_entry(0, 0, 1644, 4, 128'h40200000000000000000066d9fb);
sram_add_entry(0, 0, 1648, 4, 128'h40200000000000000000010bb50);
sram_add_entry(0, 0, 1652, 4, 128'h402000000000000000000139b8e);
sram_add_entry(0, 0, 1656, 4, 128'h40200000000000000000034094f);
sram_add_entry(0, 0, 1660, 4, 128'h402000000000000000000f852df);
sram_add_entry(0, 0, 1664, 4, 128'h402000000000000000000b4b4a5);
sram_add_entry(0, 0, 1668, 4, 128'h4020000000000000000007de478);
sram_add_entry(0, 0, 1672, 4, 128'h4020000000000000000003db18f);
sram_add_entry(0, 0, 1676, 4, 128'h402000000000000000000d272a2);
sram_add_entry(0, 0, 1680, 4, 128'h4020000000000000000008fb4b5);
sram_add_entry(0, 0, 1684, 4, 128'h40200000000000000000039e1a2);
sram_add_entry(0, 0, 1688, 4, 128'h402000000000000000000bcc07b);
sram_add_entry(0, 0, 1692, 4, 128'h402000000000000000000b2ab05);
sram_add_entry(0, 0, 1696, 4, 128'h402000000000000000000f3b478);
sram_add_entry(0, 0, 1700, 4, 128'h4020000000000000000009c9331);
sram_add_entry(0, 0, 1704, 4, 128'h4020000000000000000000570f8);
sram_add_entry(0, 0, 1708, 4, 128'h40200000000000000000092489c);
sram_add_entry(0, 0, 1712, 4, 128'h402000000000000000000d0fc4d);
sram_add_entry(0, 0, 1716, 4, 128'h4020000000000000000002acd7b);
sram_add_entry(0, 0, 1720, 4, 128'h402000000000000000000ab42dd);
sram_add_entry(0, 0, 1724, 4, 128'h402000000000000000000e77e1b);
sram_add_entry(0, 0, 1728, 4, 128'h40200000000000000000081a3c5);
sram_add_entry(0, 0, 1732, 4, 128'h4020000000000000000006cf1fa);
sram_add_entry(0, 0, 1736, 4, 128'h40200000000000000000034d05e);
sram_add_entry(0, 0, 1740, 4, 128'h4020000000000000000002b443d);
sram_add_entry(0, 0, 1744, 4, 128'h40200000000000000000097d73f);
sram_add_entry(0, 0, 1748, 4, 128'h402000000000000000000158478);
sram_add_entry(0, 0, 1752, 4, 128'h402000000000000000000e145aa);
sram_add_entry(0, 0, 1756, 4, 128'h4020000000000000000001c385e);
sram_add_entry(0, 0, 1760, 4, 128'h402000000000000000000adbce3);
sram_add_entry(0, 0, 1764, 4, 128'h402000000000000000000d72c20);
sram_add_entry(0, 0, 1768, 4, 128'h4020000000000000000005a3b1b);
sram_add_entry(0, 0, 1772, 4, 128'h4020000000000000000005eaede);
sram_add_entry(0, 0, 1776, 4, 128'h402000000000000000000651848);
sram_add_entry(0, 0, 1780, 4, 128'h402000000000000000000977b39);
sram_add_entry(0, 0, 1784, 4, 128'h4020000000000000000005cea8e);
sram_add_entry(0, 0, 1788, 4, 128'h4020000000000000000003b6c9a);
sram_add_entry(0, 0, 1792, 4, 128'h402000000000000000000492ee4);
sram_add_entry(0, 0, 1796, 4, 128'h4020000000000000000009a047c);
sram_add_entry(0, 0, 1800, 4, 128'h402000000000000000000608036);
sram_add_entry(0, 0, 1804, 4, 128'h402000000000000000000cbe70e);
sram_add_entry(0, 0, 1808, 4, 128'h4020000000000000000001eb27a);
sram_add_entry(0, 0, 1812, 4, 128'h402000000000000000000751c3a);
sram_add_entry(0, 0, 1816, 4, 128'h4020000000000000000002b749f);
sram_add_entry(0, 0, 1820, 4, 128'h4020000000000000000007ab9cd);
sram_add_entry(0, 0, 1824, 4, 128'h402000000000000000000db74b0);
sram_add_entry(0, 0, 1828, 4, 128'h40200000000000000000038ccf5);
sram_add_entry(0, 0, 1832, 4, 128'h402000000000000000000b81901);
sram_add_entry(0, 0, 1836, 4, 128'h402000000000000000000db6f8a);
sram_add_entry(0, 0, 1840, 4, 128'h402000000000000000000bdfaee);
sram_add_entry(0, 0, 1844, 4, 128'h402000000000000000000ab9134);
sram_add_entry(0, 0, 1848, 4, 128'h4020000000000000000006d74aa);
sram_add_entry(0, 0, 1852, 4, 128'h402000000000000000000f71076);
sram_add_entry(0, 0, 1856, 4, 128'h402000000000000000000579bdc);
sram_add_entry(0, 0, 1860, 4, 128'h402000000000000000000bbbd64);
sram_add_entry(0, 0, 1864, 4, 128'h40200000000000000000083ae74);
sram_add_entry(0, 0, 1868, 4, 128'h402000000000000000000f8c1d9);
sram_add_entry(0, 0, 1872, 4, 128'h402000000000000000000c8ed3e);
sram_add_entry(0, 0, 1876, 4, 128'h4020000000000000000002bf8dc);
sram_add_entry(0, 0, 1880, 4, 128'h40200000000000000000016e5de);
sram_add_entry(0, 0, 1884, 4, 128'h402000000000000000000b99492);
sram_add_entry(0, 0, 1888, 4, 128'h402000000000000000000820b16);
sram_add_entry(0, 0, 1892, 4, 128'h4020000000000000000008ae9cf);
sram_add_entry(0, 0, 1896, 4, 128'h402000000000000000000f6aad1);
sram_add_entry(0, 0, 1900, 4, 128'h402000000000000000000def433);
sram_add_entry(0, 0, 1904, 4, 128'h40200000000000000000060e02b);
sram_add_entry(0, 0, 1908, 4, 128'h402000000000000000000ba10d9);
sram_add_entry(0, 0, 1912, 4, 128'h402000000000000000000125ae0);
sram_add_entry(0, 0, 1916, 4, 128'h40200000000000000000075abca);
sram_add_entry(0, 0, 1920, 4, 128'h4020000000000000000007d0a37);
sram_add_entry(0, 0, 1924, 4, 128'h40200000000000000000076c3eb);
sram_add_entry(0, 0, 1928, 4, 128'h402000000000000000000ee5867);
sram_add_entry(0, 0, 1932, 4, 128'h402000000000000000000a63aa9);
sram_add_entry(0, 0, 1936, 4, 128'h4020000000000000000003bf1a7);
sram_add_entry(0, 0, 1940, 4, 128'h40200000000000000000041b00e);
sram_add_entry(0, 0, 1944, 4, 128'h4020000000000000000005dfcea);
sram_add_entry(0, 0, 1948, 4, 128'h402000000000000000000856939);
sram_add_entry(0, 0, 1952, 4, 128'h40200000000000000000007fdd0);
sram_add_entry(0, 0, 1956, 4, 128'h402000000000000000000cac855);
sram_add_entry(0, 0, 1960, 4, 128'h40200000000000000000082c86b);
sram_add_entry(0, 0, 1964, 4, 128'h4020000000000000000007d64e0);
sram_add_entry(0, 0, 1968, 4, 128'h402000000000000000000c05790);
sram_add_entry(0, 0, 1972, 4, 128'h40200000000000000000041b488);
sram_add_entry(0, 0, 1976, 4, 128'h40200000000000000000019ef12);
sram_add_entry(0, 0, 1980, 4, 128'h40200000000000000000089d14b);
sram_add_entry(0, 0, 1984, 4, 128'h402000000000000000000b42732);
sram_add_entry(0, 0, 1988, 4, 128'h402000000000000000000a795fa);
sram_add_entry(0, 0, 1992, 4, 128'h402000000000000000000a72e70);
sram_add_entry(0, 0, 1996, 4, 128'h402000000000000000000a16e73);
sram_add_entry(0, 0, 2000, 4, 128'h40200000000000000000080fe5c);
sram_add_entry(0, 0, 2004, 4, 128'h402000000000000000000bdf1f7);
sram_add_entry(0, 0, 2008, 4, 128'h40200000000000000000024e03d);
sram_add_entry(0, 0, 2012, 4, 128'h402000000000000000000cd8833);
sram_add_entry(0, 0, 2016, 4, 128'h402000000000000000000d48427);
sram_add_entry(0, 0, 2020, 4, 128'h40200000000000000000029413e);
sram_add_entry(0, 0, 2024, 4, 128'h40200000000000000000099f215);
sram_add_entry(0, 0, 2028, 4, 128'h40200000000000000000043ea2c);
sram_add_entry(0, 0, 2032, 4, 128'h402000000000000000000b05ed6);
sram_add_entry(0, 0, 2036, 4, 128'h402000000000000000000359c4e);
sram_add_entry(0, 0, 2040, 4, 128'h402000000000000000000a53a50);
sram_add_entry(0, 0, 2044, 4, 128'h402000000000000000000ba0217);
sram_add_entry(0, 0, 2048, 4, 128'h402000000000000000000a7a8be);
sram_add_entry(0, 0, 2052, 4, 128'h402000000000000000000117261);
sram_add_entry(0, 0, 2056, 4, 128'h402000000000000000000ba40b1);
sram_add_entry(0, 0, 2060, 4, 128'h402000000000000000000d3778c);
sram_add_entry(0, 0, 2064, 4, 128'h402000000000000000000133300);
sram_add_entry(0, 0, 2068, 4, 128'h4020000000000000000008026d0);
sram_add_entry(0, 0, 2072, 4, 128'h4020000000000000000003c2a96);
sram_add_entry(0, 0, 2076, 4, 128'h402000000000000000000af2172);
sram_add_entry(0, 0, 2080, 4, 128'h402000000000000000000f83e69);
sram_add_entry(0, 0, 2084, 4, 128'h4020000000000000000002bae72);
sram_add_entry(0, 0, 2088, 4, 128'h402000000000000000000aaffe3);
sram_add_entry(0, 0, 2092, 4, 128'h402000000000000000000e47a3a);
sram_add_entry(0, 0, 2096, 4, 128'h402000000000000000000ecf185);
sram_add_entry(0, 0, 2100, 4, 128'h4020000000000000000002ed0f5);
sram_add_entry(0, 0, 2104, 4, 128'h402000000000000000000d53425);
sram_add_entry(0, 0, 2108, 4, 128'h402000000000000000000ecfd2a);
sram_add_entry(0, 0, 2112, 4, 128'h402000000000000000000c133a2);
sram_add_entry(0, 0, 2116, 4, 128'h402000000000000000000b51947);
sram_add_entry(0, 0, 2120, 4, 128'h4020000000000000000001f5b10);
sram_add_entry(0, 0, 2124, 4, 128'h402000000000000000000724175);
sram_add_entry(0, 0, 2128, 4, 128'h4020000000000000000004a6946);
sram_add_entry(0, 0, 2132, 4, 128'h402000000000000000000f4634a);
sram_add_entry(0, 0, 2136, 4, 128'h40200000000000000000074e5f6);
sram_add_entry(0, 0, 2140, 4, 128'h402000000000000000000b53980);
sram_add_entry(0, 0, 2144, 4, 128'h402000000000000000000bbd32a);
sram_add_entry(0, 0, 2148, 4, 128'h4020000000000000000004beff2);
sram_add_entry(0, 0, 2152, 4, 128'h402000000000000000000c8358f);
sram_add_entry(0, 0, 2156, 4, 128'h402000000000000000000cb9cd4);
sram_add_entry(0, 0, 2160, 4, 128'h4020000000000000000005a3371);
sram_add_entry(0, 0, 2164, 4, 128'h402000000000000000000b24300);
sram_add_entry(0, 0, 2168, 4, 128'h4020000000000000000001fb996);
sram_add_entry(0, 0, 2172, 4, 128'h402000000000000000000bd4f61);
sram_add_entry(0, 0, 2176, 4, 128'h4020000000000000000008abbcd);
sram_add_entry(0, 0, 2180, 4, 128'h402000000000000000000b9b2c6);
sram_add_entry(0, 0, 2184, 4, 128'h402000000000000000000638408);
sram_add_entry(0, 0, 2188, 4, 128'h402000000000000000000d821e0);
sram_add_entry(0, 0, 2192, 4, 128'h402000000000000000000694d89);
sram_add_entry(0, 0, 2196, 4, 128'h402000000000000000000cc2430);
sram_add_entry(0, 0, 2200, 4, 128'h4020000000000000000000b3c95);
sram_add_entry(0, 0, 2204, 4, 128'h4020000000000000000002c40c9);
sram_add_entry(0, 0, 2208, 4, 128'h402000000000000000000ec7053);
sram_add_entry(0, 0, 2212, 4, 128'h4020000000000000000008adfbd);
sram_add_entry(0, 0, 2216, 4, 128'h40200000000000000000015e421);
sram_add_entry(0, 0, 2220, 4, 128'h402000000000000000000cd639d);
sram_add_entry(0, 0, 2224, 4, 128'h40200000000000000000006a5ec);
sram_add_entry(0, 0, 2228, 4, 128'h4020000000000000000004837b3);
sram_add_entry(0, 0, 2232, 4, 128'h4020000000000000000003c1296);
sram_add_entry(0, 0, 2236, 4, 128'h4020000000000000000009854db);
sram_add_entry(0, 0, 2240, 4, 128'h402000000000000000000e23953);
sram_add_entry(0, 0, 2244, 4, 128'h4020000000000000000006e5f61);
sram_add_entry(0, 0, 2248, 4, 128'h402000000000000000000b67704);
sram_add_entry(0, 0, 2252, 4, 128'h402000000000000000000c188f5);
sram_add_entry(0, 0, 2256, 4, 128'h4020000000000000000009f0af0);
sram_add_entry(0, 0, 2260, 4, 128'h40200000000000000000013deba);
sram_add_entry(0, 0, 2264, 4, 128'h402000000000000000000d836a2);
sram_add_entry(0, 0, 2268, 4, 128'h402000000000000000000378015);
sram_add_entry(0, 0, 2272, 4, 128'h40200000000000000000006857c);
sram_add_entry(0, 0, 2276, 4, 128'h402000000000000000000920848);
sram_add_entry(0, 0, 2280, 4, 128'h402000000000000000000df91e5);
sram_add_entry(0, 0, 2284, 4, 128'h402000000000000000000203539);
sram_add_entry(0, 0, 2288, 4, 128'h402000000000000000000e0e16e);
sram_add_entry(0, 0, 2292, 4, 128'h402000000000000000000518348);
sram_add_entry(0, 0, 2296, 4, 128'h40200000000000000000029589f);
sram_add_entry(0, 0, 2300, 4, 128'h402000000000000000000d5eff5);
sram_add_entry(0, 0, 2304, 4, 128'h402000000000000000000a8909a);
sram_add_entry(0, 0, 2308, 4, 128'h402000000000000000000c6ccb7);
sram_add_entry(0, 0, 2312, 4, 128'h4020000000000000000008fd56d);
sram_add_entry(0, 0, 2316, 4, 128'h402000000000000000000bf7f6d);
sram_add_entry(0, 0, 2320, 4, 128'h4020000000000000000006a229b);
sram_add_entry(0, 0, 2324, 4, 128'h402000000000000000000a7dd84);
sram_add_entry(0, 0, 2328, 4, 128'h4020000000000000000003d9854);
sram_add_entry(0, 0, 2332, 4, 128'h4020000000000000000003c87c6);
sram_add_entry(0, 0, 2336, 4, 128'h402000000000000000000588ad5);
sram_add_entry(0, 0, 2340, 4, 128'h402000000000000000000eaaf14);
sram_add_entry(0, 0, 2344, 4, 128'h402000000000000000000344bf2);
sram_add_entry(0, 0, 2348, 4, 128'h4020000000000000000003d9161);
sram_add_entry(0, 0, 2352, 4, 128'h4020000000000000000000415ce);
sram_add_entry(0, 0, 2356, 4, 128'h4020000000000000000000b69cc);
sram_add_entry(0, 0, 2360, 4, 128'h402000000000000000000fe9312);
sram_add_entry(0, 0, 2364, 4, 128'h402000000000000000000878cb6);
sram_add_entry(0, 0, 2368, 4, 128'h40200000000000000000038cf4e);
sram_add_entry(0, 0, 2372, 4, 128'h40200000000000000000076dcb4);
sram_add_entry(0, 0, 2376, 4, 128'h402000000000000000000702f85);
sram_add_entry(0, 0, 2380, 4, 128'h402000000000000000000ecdc20);
sram_add_entry(0, 0, 2384, 4, 128'h402000000000000000000064eed);
sram_add_entry(0, 0, 2388, 4, 128'h402000000000000000000197ad7);
sram_add_entry(0, 0, 2392, 4, 128'h402000000000000000000860fe2);
sram_add_entry(0, 0, 2396, 4, 128'h402000000000000000000aafcfa);
sram_add_entry(0, 0, 2400, 4, 128'h402000000000000000000b3fdf0);
sram_add_entry(0, 0, 2404, 4, 128'h402000000000000000000075513);
sram_add_entry(0, 0, 2408, 4, 128'h40200000000000000000013141b);
sram_add_entry(0, 0, 2412, 4, 128'h402000000000000000000d07c80);
sram_add_entry(0, 0, 2416, 4, 128'h4020000000000000000007023d5);
sram_add_entry(0, 0, 2420, 4, 128'h40200000000000000000088bbc7);
sram_add_entry(0, 0, 2424, 4, 128'h4020000000000000000008bd1c2);
sram_add_entry(0, 0, 2428, 4, 128'h402000000000000000000ede0cc);
sram_add_entry(0, 0, 2432, 4, 128'h40200000000000000000011d1b8);
sram_add_entry(0, 0, 2436, 4, 128'h402000000000000000000d0feb3);
sram_add_entry(0, 0, 2440, 4, 128'h402000000000000000000ef7aab);
sram_add_entry(0, 0, 2444, 4, 128'h402000000000000000000929846);
sram_add_entry(0, 0, 2448, 4, 128'h40200000000000000000087f8f5);
sram_add_entry(0, 0, 2452, 4, 128'h402000000000000000000f6d906);
sram_add_entry(0, 0, 2456, 4, 128'h402000000000000000000301023);
sram_add_entry(0, 0, 2460, 4, 128'h402000000000000000000c0367e);
sram_add_entry(0, 0, 2464, 4, 128'h4020000000000000000000b5225);
sram_add_entry(0, 0, 2468, 4, 128'h4020000000000000000001abda8);
sram_add_entry(0, 0, 2472, 4, 128'h402000000000000000000f76cf7);
sram_add_entry(0, 0, 2476, 4, 128'h402000000000000000000715672);
sram_add_entry(0, 0, 2480, 4, 128'h4020000000000000000007a6132);
sram_add_entry(0, 0, 2484, 4, 128'h402000000000000000000443d93);
sram_add_entry(0, 0, 2488, 4, 128'h402000000000000000000eb213b);
sram_add_entry(0, 0, 2492, 4, 128'h4020000000000000000004d47a0);
sram_add_entry(0, 0, 2496, 4, 128'h402000000000000000000a05377);
sram_add_entry(0, 0, 2500, 4, 128'h4020000000000000000006ac1b8);
sram_add_entry(0, 0, 2504, 4, 128'h4020000000000000000007a773d);
sram_add_entry(0, 0, 2508, 4, 128'h402000000000000000000e5e3a5);
sram_add_entry(0, 0, 2512, 4, 128'h402000000000000000000c9746b);
sram_add_entry(0, 0, 2516, 4, 128'h40200000000000000000023a9d3);
sram_add_entry(0, 0, 2520, 4, 128'h4020000000000000000004ec356);
sram_add_entry(0, 0, 2524, 4, 128'h402000000000000000000075d68);
sram_add_entry(0, 0, 2528, 4, 128'h4020000000000000000003f8eba);
sram_add_entry(0, 0, 2532, 4, 128'h4020000000000000000004d98e8);
sram_add_entry(0, 0, 2536, 4, 128'h40200000000000000000098da92);
sram_add_entry(0, 0, 2540, 4, 128'h402000000000000000000ca02ef);
sram_add_entry(0, 0, 2544, 4, 128'h402000000000000000000924656);
sram_add_entry(0, 0, 2548, 4, 128'h4020000000000000000004eb306);
sram_add_entry(0, 0, 2552, 4, 128'h40200000000000000000033a608);
sram_add_entry(0, 0, 2556, 4, 128'h402000000000000000000291e21);
sram_add_entry(0, 0, 2560, 4, 128'h402000000000000000000c4dc56);
sram_add_entry(0, 0, 2564, 4, 128'h4020000000000000000001b53a4);
sram_add_entry(0, 0, 2568, 4, 128'h40200000000000000000009d22f);
sram_add_entry(0, 0, 2572, 4, 128'h4020000000000000000005a1b8f);
sram_add_entry(0, 0, 2576, 4, 128'h402000000000000000000e01679);
sram_add_entry(0, 0, 2580, 4, 128'h40200000000000000000044e0ed);
sram_add_entry(0, 0, 2584, 4, 128'h402000000000000000000c9bb74);
sram_add_entry(0, 0, 2588, 4, 128'h4020000000000000000005c1683);
sram_add_entry(0, 0, 2592, 4, 128'h4020000000000000000005fbc9d);
sram_add_entry(0, 0, 2596, 4, 128'h402000000000000000000bc2b03);
sram_add_entry(0, 0, 2600, 4, 128'h40200000000000000000044df86);
sram_add_entry(0, 0, 2604, 4, 128'h402000000000000000000dadec5);
sram_add_entry(0, 0, 2608, 4, 128'h4020000000000000000002fa3c2);
sram_add_entry(0, 0, 2612, 4, 128'h402000000000000000000795c0b);
sram_add_entry(0, 0, 2616, 4, 128'h402000000000000000000c6f84e);
sram_add_entry(0, 0, 2620, 4, 128'h402000000000000000000b16934);
sram_add_entry(0, 0, 2624, 4, 128'h4020000000000000000009460ec);
sram_add_entry(0, 0, 2628, 4, 128'h402000000000000000000961e88);
sram_add_entry(0, 0, 2632, 4, 128'h402000000000000000000c93603);
sram_add_entry(0, 0, 2636, 4, 128'h402000000000000000000f71bb0);
sram_add_entry(0, 0, 2640, 4, 128'h402000000000000000000b1611c);
sram_add_entry(0, 0, 2644, 4, 128'h402000000000000000000ec7932);
sram_add_entry(0, 0, 2648, 4, 128'h40200000000000000000043bb09);
sram_add_entry(0, 0, 2652, 4, 128'h402000000000000000000040cb8);
sram_add_entry(0, 0, 2656, 4, 128'h40200000000000000000085d475);
sram_add_entry(0, 0, 2660, 4, 128'h402000000000000000000a661a8);
sram_add_entry(0, 0, 2664, 4, 128'h4020000000000000000000f38b5);
sram_add_entry(0, 0, 2668, 4, 128'h402000000000000000000986622);
sram_add_entry(0, 0, 2672, 4, 128'h40200000000000000000072876e);
sram_add_entry(0, 0, 2676, 4, 128'h40200000000000000000026c981);
sram_add_entry(0, 0, 2680, 4, 128'h402000000000000000000c3c23a);
sram_add_entry(0, 0, 2684, 4, 128'h402000000000000000000907259);
sram_add_entry(0, 0, 2688, 4, 128'h40200000000000000000052165d);
sram_add_entry(0, 0, 2692, 4, 128'h40200000000000000000095fcd7);
sram_add_entry(0, 0, 2696, 4, 128'h4020000000000000000002dc5de);
sram_add_entry(0, 0, 2700, 4, 128'h4020000000000000000003bd5a3);
sram_add_entry(0, 0, 2704, 4, 128'h402000000000000000000a551ba);
sram_add_entry(0, 0, 2708, 4, 128'h40200000000000000000035e5cb);
sram_add_entry(0, 0, 2712, 4, 128'h402000000000000000000c960bd);
sram_add_entry(0, 0, 2716, 4, 128'h40200000000000000000023b8b6);
sram_add_entry(0, 0, 2720, 4, 128'h402000000000000000000d4d778);
sram_add_entry(0, 0, 2724, 4, 128'h402000000000000000000ea3ee3);
sram_add_entry(0, 0, 2728, 4, 128'h4020000000000000000001d84d3);
sram_add_entry(0, 0, 2732, 4, 128'h40200000000000000000077135c);
sram_add_entry(0, 0, 2736, 4, 128'h40200000000000000000061df00);
sram_add_entry(0, 0, 2740, 4, 128'h402000000000000000000a9a5bc);
sram_add_entry(0, 0, 2744, 4, 128'h402000000000000000000ba4d19);
sram_add_entry(0, 0, 2748, 4, 128'h402000000000000000000ccf409);
sram_add_entry(0, 0, 2752, 4, 128'h40200000000000000000085da8d);
sram_add_entry(0, 0, 2756, 4, 128'h402000000000000000000615d80);
sram_add_entry(0, 0, 2760, 4, 128'h402000000000000000000726469);
sram_add_entry(0, 0, 2764, 4, 128'h40200000000000000000069cc0a);
sram_add_entry(0, 0, 2768, 4, 128'h402000000000000000000b23db7);
sram_add_entry(0, 0, 2772, 4, 128'h402000000000000000000512c45);
sram_add_entry(0, 0, 2776, 4, 128'h402000000000000000000dcffc3);
sram_add_entry(0, 0, 2780, 4, 128'h402000000000000000000cc8fd4);
sram_add_entry(0, 0, 2784, 4, 128'h402000000000000000000ac910e);
sram_add_entry(0, 0, 2788, 4, 128'h40200000000000000000066efed);
sram_add_entry(0, 0, 2792, 4, 128'h402000000000000000000d0094e);
sram_add_entry(0, 0, 2796, 4, 128'h402000000000000000000c23370);
sram_add_entry(0, 0, 2800, 4, 128'h402000000000000000000ace597);
sram_add_entry(0, 3, 0, 4, 128'h7ab000000000000000000deadbf);
sram_add_entry(0, 3, 4, 4, 128'h4030000000000000000b54f67e3);
sram_add_entry(0, 3, 8, 4, 128'h403000000000000000082701ad9);
sram_add_entry(0, 3, 12, 4, 128'h403000000000000000073a0f3c7);
sram_add_entry(0, 3, 16, 4, 128'h4030000000000000000094c7976);
sram_add_entry(0, 3, 20, 4, 128'h4030000000000000000ce105c36);
sram_add_entry(0, 3, 24, 4, 128'h4030000000000000000b834579a);
sram_add_entry(0, 3, 28, 4, 128'h40300000000000000006b75275d);
sram_add_entry(0, 3, 32, 4, 128'h403000000000000000065729ff2);
sram_add_entry(0, 3, 36, 4, 128'h403000000000000000009c97d69);
sram_add_entry(0, 3, 40, 4, 128'h403000000000000000095f0765a);
sram_add_entry(0, 3, 44, 4, 128'h4030000000000000000c6cb3d40);
sram_add_entry(0, 3, 48, 4, 128'h403000000000000000051099d25);
sram_add_entry(0, 3, 52, 4, 128'h403000000000000000013be202f);
sram_add_entry(0, 3, 56, 4, 128'h4030000000000000000aded021e);
sram_add_entry(0, 3, 60, 4, 128'h4030000000000000000a8ab1332);
sram_add_entry(0, 3, 64, 4, 128'h4030000000000000000dee9be17);
sram_add_entry(0, 3, 68, 4, 128'h403000000000000000010344d26);
sram_add_entry(0, 3, 72, 4, 128'h4030000000000000000eee66d45);
sram_add_entry(0, 3, 76, 4, 128'h403000000000000000085015a63);
sram_add_entry(0, 3, 80, 4, 128'h403000000000000000011b09ad8);
sram_add_entry(0, 3, 84, 4, 128'h403000000000000000095ed2ba2);
sram_add_entry(0, 3, 88, 4, 128'h4030000000000000000ae60dfc5);
sram_add_entry(0, 3, 92, 4, 128'h4030000000000000000f32db0c1);
sram_add_entry(0, 3, 96, 4, 128'h40300000000000000009d50520d);
sram_add_entry(0, 3, 100, 4, 128'h403000000000000000083fa86a3);
sram_add_entry(0, 3, 104, 4, 128'h4030000000000000000fed13352);
sram_add_entry(0, 3, 108, 4, 128'h40300000000000000006c4cf1a3);
sram_add_entry(0, 3, 112, 4, 128'h40300000000000000001e12a2c3);
sram_add_entry(0, 3, 116, 4, 128'h4030000000000000000b199f9bd);
sram_add_entry(0, 3, 120, 4, 128'h40300000000000000005edff01d);
sram_add_entry(0, 3, 124, 4, 128'h4030000000000000000777705d7);
sram_add_entry(0, 3, 128, 4, 128'h403000000000000000065c1fcdf);
sram_add_entry(0, 3, 132, 4, 128'h403000000000000000037860217);
sram_add_entry(0, 3, 136, 4, 128'h403000000000000000060b3521a);
sram_add_entry(0, 3, 140, 4, 128'h40300000000000000000d2e417a);
sram_add_entry(0, 3, 144, 4, 128'h40300000000000000000e4f4fa6);
sram_add_entry(0, 3, 148, 4, 128'h403000000000000000056ca43a2);
sram_add_entry(0, 3, 152, 4, 128'h4030000000000000000a3d16cc5);
sram_add_entry(0, 3, 156, 4, 128'h403000000000000000017fdfddb);
sram_add_entry(0, 3, 160, 4, 128'h40300000000000000008dc5fc1e);
sram_add_entry(0, 3, 164, 4, 128'h4030000000000000000dda06a7d);
sram_add_entry(0, 3, 168, 4, 128'h4030000000000000000ee1abcfe);
sram_add_entry(0, 3, 172, 4, 128'h4030000000000000000b6b2c311);
sram_add_entry(0, 3, 176, 4, 128'h40300000000000000005222e309);
sram_add_entry(0, 3, 180, 4, 128'h40300000000000000004de83400);
sram_add_entry(0, 3, 184, 4, 128'h4030000000000000000f55ce23a);
sram_add_entry(0, 3, 188, 4, 128'h4030000000000000000923f30a1);
sram_add_entry(0, 3, 192, 4, 128'h403000000000000000002805970);
sram_add_entry(0, 3, 196, 4, 128'h4030000000000000000600e6cd3);
sram_add_entry(0, 3, 200, 4, 128'h4030000000000000000560660db);
sram_add_entry(0, 3, 204, 4, 128'h4030000000000000000e78a38a2);
sram_add_entry(0, 3, 208, 4, 128'h4030000000000000000a2af2509);
sram_add_entry(0, 3, 212, 4, 128'h4030000000000000000bce83038);
sram_add_entry(0, 3, 216, 4, 128'h4030000000000000000c6c499c6);
sram_add_entry(0, 3, 220, 4, 128'h4030000000000000000cfe4fdb8);
sram_add_entry(0, 3, 224, 4, 128'h4030000000000000000e84582e1);
sram_add_entry(0, 3, 228, 4, 128'h40300000000000000001cbd8994);
sram_add_entry(0, 3, 232, 4, 128'h40300000000000000008725b8fe);
sram_add_entry(0, 3, 236, 4, 128'h4030000000000000000820f2dae);
sram_add_entry(0, 3, 240, 4, 128'h4030000000000000000b9ebe16e);
sram_add_entry(0, 3, 244, 4, 128'h40300000000000000008f276dcf);
sram_add_entry(0, 3, 248, 4, 128'h40300000000000000008158b691);
sram_add_entry(0, 3, 252, 4, 128'h4030000000000000000f40e5df3);
sram_add_entry(0, 3, 256, 4, 128'h40300000000000000007f3fd2ce);
sram_add_entry(0, 3, 260, 4, 128'h4030000000000000000fb50a4cb);
sram_add_entry(0, 3, 264, 4, 128'h4030000000000000000a23f290a);
sram_add_entry(0, 3, 268, 4, 128'h4030000000000000000a249d8fe);
sram_add_entry(0, 3, 272, 4, 128'h403000000000000000073ddd4d9);
sram_add_entry(0, 3, 276, 4, 128'h40300000000000000003d4518bb);
sram_add_entry(0, 3, 280, 4, 128'h4030000000000000000b12418a1);
sram_add_entry(0, 3, 284, 4, 128'h40300000000000000002b0255f5);
sram_add_entry(0, 3, 288, 4, 128'h4030000000000000000b26dbe7a);
sram_add_entry(0, 3, 292, 4, 128'h4030000000000000000be63e546);
sram_add_entry(0, 3, 296, 4, 128'h4030000000000000000ced8a116);
sram_add_entry(0, 3, 300, 4, 128'h4030000000000000000d4fd6330);
sram_add_entry(0, 3, 304, 4, 128'h403000000000000000089538b5c);
sram_add_entry(0, 3, 308, 4, 128'h40300000000000000007545692b);
sram_add_entry(0, 3, 312, 4, 128'h40300000000000000006e3d0ccd);
sram_add_entry(0, 3, 316, 4, 128'h40300000000000000001f95de86);
sram_add_entry(0, 3, 320, 4, 128'h403000000000000000032b5bb45);
sram_add_entry(0, 3, 324, 4, 128'h4030000000000000000f78ec26e);
sram_add_entry(0, 3, 328, 4, 128'h40300000000000000006a4b0fd1);
sram_add_entry(0, 3, 332, 4, 128'h40300000000000000001cb2bf20);
sram_add_entry(0, 3, 336, 4, 128'h4030000000000000000ba9bed68);
sram_add_entry(0, 3, 340, 4, 128'h4030000000000000000a559577e);
sram_add_entry(0, 3, 344, 4, 128'h403000000000000000090bad641);
sram_add_entry(0, 3, 348, 4, 128'h4030000000000000000f6c3245a);
sram_add_entry(0, 3, 352, 4, 128'h4030000000000000000ecda72aa);
sram_add_entry(0, 3, 356, 4, 128'h4030000000000000000b3b7c2b4);
sram_add_entry(0, 3, 360, 4, 128'h40300000000000000001428e333);
sram_add_entry(0, 3, 364, 4, 128'h40300000000000000005b902d27);
sram_add_entry(0, 3, 368, 4, 128'h4030000000000000000153d8c14);
sram_add_entry(0, 3, 372, 4, 128'h403000000000000000092d06347);
sram_add_entry(0, 3, 376, 4, 128'h40300000000000000002c2c4397);
sram_add_entry(0, 3, 380, 4, 128'h4030000000000000000b7423e69);
sram_add_entry(0, 3, 384, 4, 128'h4030000000000000000015a6481);
sram_add_entry(0, 3, 388, 4, 128'h4030000000000000000dfb988cd);
sram_add_entry(0, 3, 392, 4, 128'h4030000000000000000cde361c7);
sram_add_entry(0, 3, 396, 4, 128'h4030000000000000000e308f937);
sram_add_entry(0, 3, 400, 4, 128'h40300000000000000002164ee50);
sram_add_entry(0, 3, 404, 4, 128'h4030000000000000000616c5a7f);
sram_add_entry(0, 3, 408, 4, 128'h4030000000000000000db1b964e);
sram_add_entry(0, 3, 412, 4, 128'h40300000000000000005154a7da);
sram_add_entry(0, 3, 416, 4, 128'h40300000000000000005c6ec2c4);
sram_add_entry(0, 3, 420, 4, 128'h40300000000000000004294e76d);
sram_add_entry(0, 3, 424, 4, 128'h40300000000000000005220f2ca);
sram_add_entry(0, 3, 428, 4, 128'h4030000000000000000da566993);
sram_add_entry(0, 3, 432, 4, 128'h40300000000000000001d318de4);
sram_add_entry(0, 3, 436, 4, 128'h40300000000000000003346495f);
sram_add_entry(0, 3, 440, 4, 128'h4030000000000000000f4a6db31);
sram_add_entry(0, 3, 444, 4, 128'h40300000000000000001e9b4645);
sram_add_entry(0, 3, 448, 4, 128'h4030000000000000000c1ce109e);
sram_add_entry(0, 3, 452, 4, 128'h403000000000000000093229de8);
sram_add_entry(0, 3, 456, 4, 128'h403000000000000000011553172);
sram_add_entry(0, 3, 460, 4, 128'h40300000000000000005db88c38);
sram_add_entry(0, 3, 464, 4, 128'h40300000000000000002968364c);
sram_add_entry(0, 3, 468, 4, 128'h40300000000000000009c14bafb);
sram_add_entry(0, 3, 472, 4, 128'h4030000000000000000115ed45f);
sram_add_entry(0, 3, 476, 4, 128'h4030000000000000000c528fcec);
sram_add_entry(0, 3, 480, 4, 128'h40300000000000000002ea562ca);
sram_add_entry(0, 3, 484, 4, 128'h403000000000000000070397c26);
sram_add_entry(0, 3, 488, 4, 128'h403000000000000000017516503);
sram_add_entry(0, 3, 492, 4, 128'h4030000000000000000e2648a6b);
sram_add_entry(0, 3, 496, 4, 128'h40300000000000000009050a552);
sram_add_entry(0, 3, 500, 4, 128'h40300000000000000002ae6316d);
sram_add_entry(0, 3, 504, 4, 128'h403000000000000000085b27335);
sram_add_entry(0, 3, 508, 4, 128'h4030000000000000000edcea4e9);
sram_add_entry(0, 3, 512, 4, 128'h4030000000000000000c3666129);
sram_add_entry(0, 3, 516, 4, 128'h4030000000000000000dde557c9);
sram_add_entry(0, 3, 520, 4, 128'h403000000000000000036fcd376);
sram_add_entry(0, 3, 524, 4, 128'h4030000000000000000d0642c0d);
sram_add_entry(0, 3, 528, 4, 128'h40300000000000000005191ba09);
sram_add_entry(0, 3, 532, 4, 128'h4030000000000000000307e4946);
sram_add_entry(0, 3, 536, 4, 128'h403000000000000000041821824);
sram_add_entry(0, 3, 540, 4, 128'h4030000000000000000787c80c6);
sram_add_entry(0, 3, 544, 4, 128'h4030000000000000000f618f71d);
sram_add_entry(0, 3, 548, 4, 128'h4030000000000000000edacc3d3);
sram_add_entry(0, 3, 552, 4, 128'h40300000000000000007e52d942);
sram_add_entry(0, 3, 556, 4, 128'h40300000000000000003f71fbaf);
sram_add_entry(0, 3, 560, 4, 128'h403000000000000000023350757);
sram_add_entry(0, 3, 564, 4, 128'h4030000000000000000652439de);
sram_add_entry(0, 3, 568, 4, 128'h403000000000000000067c671d1);
sram_add_entry(0, 3, 572, 4, 128'h403000000000000000059998fe8);
sram_add_entry(0, 3, 576, 4, 128'h4030000000000000000d3f88f1f);
sram_add_entry(0, 3, 580, 4, 128'h4030000000000000000c2b4ab74);
sram_add_entry(0, 3, 584, 4, 128'h4030000000000000000abc85eb1);
sram_add_entry(0, 3, 588, 4, 128'h4030000000000000000464a1392);
sram_add_entry(0, 3, 592, 4, 128'h403000000000000000091c8a041);
sram_add_entry(0, 3, 596, 4, 128'h40300000000000000008224a2e1);
sram_add_entry(0, 3, 600, 4, 128'h4030000000000000000e4590888);
sram_add_entry(0, 3, 604, 4, 128'h4030000000000000000ec9ac7c1);
sram_add_entry(0, 3, 608, 4, 128'h403000000000000000066424878);
sram_add_entry(0, 3, 612, 4, 128'h403000000000000000067af253d);
sram_add_entry(0, 3, 616, 4, 128'h403000000000000000045d5dbde);
sram_add_entry(0, 3, 620, 4, 128'h4030000000000000000c54a488a);
sram_add_entry(0, 3, 624, 4, 128'h4030000000000000000ee973819);
sram_add_entry(0, 3, 628, 4, 128'h4030000000000000000f58cfd37);
sram_add_entry(0, 3, 632, 4, 128'h4030000000000000000574bcdc4);
sram_add_entry(0, 3, 636, 4, 128'h4030000000000000000a7a8595a);
sram_add_entry(0, 3, 640, 4, 128'h4030000000000000000d3b139e9);
sram_add_entry(0, 3, 644, 4, 128'h40300000000000000006e36b346);
sram_add_entry(0, 3, 648, 4, 128'h4030000000000000000da8acfb4);
sram_add_entry(0, 3, 652, 4, 128'h4030000000000000000185f3089);
sram_add_entry(0, 3, 656, 4, 128'h4030000000000000000bde907e3);
sram_add_entry(0, 3, 660, 4, 128'h403000000000000000004d5fbad);
sram_add_entry(0, 3, 664, 4, 128'h4030000000000000000ab507ea2);
sram_add_entry(0, 3, 668, 4, 128'h40300000000000000006e8feba1);
sram_add_entry(0, 3, 672, 4, 128'h4030000000000000000d2a5d8f4);
sram_add_entry(0, 3, 676, 4, 128'h40300000000000000001f98cf7f);
sram_add_entry(0, 3, 680, 4, 128'h4030000000000000000e00933b5);
sram_add_entry(0, 3, 684, 4, 128'h403000000000000000094318208);
sram_add_entry(0, 3, 688, 4, 128'h40300000000000000005eef8c5a);
sram_add_entry(0, 3, 692, 4, 128'h4030000000000000000fb9a2b06);
sram_add_entry(0, 3, 696, 4, 128'h40300000000000000001dbc0c13);
sram_add_entry(0, 3, 700, 4, 128'h403000000000000000096e2cec1);
sram_add_entry(0, 3, 704, 4, 128'h4030000000000000000bbfa2397);
sram_add_entry(0, 3, 708, 4, 128'h40300000000000000001284be5f);
sram_add_entry(0, 3, 712, 4, 128'h4030000000000000000b20a2de4);
sram_add_entry(0, 3, 716, 4, 128'h4030000000000000000521ee751);
sram_add_entry(0, 3, 720, 4, 128'h403000000000000000084d1e904);
sram_add_entry(0, 3, 724, 4, 128'h4030000000000000000be957768);
sram_add_entry(0, 3, 728, 4, 128'h403000000000000000083a7c5dc);
sram_add_entry(0, 3, 732, 4, 128'h40300000000000000005ef8ecda);
sram_add_entry(0, 3, 736, 4, 128'h4030000000000000000c9ef88d4);
sram_add_entry(0, 3, 740, 4, 128'h4030000000000000000dba7c009);
sram_add_entry(0, 3, 744, 4, 128'h40300000000000000006a4242f9);
sram_add_entry(0, 3, 748, 4, 128'h4030000000000000000cb1f7db1);
sram_add_entry(0, 3, 752, 4, 128'h4030000000000000000282df15a);
sram_add_entry(0, 3, 756, 4, 128'h403000000000000000011da4159);
sram_add_entry(0, 3, 760, 4, 128'h4030000000000000000c979d2c0);
sram_add_entry(0, 3, 764, 4, 128'h403000000000000000015d0a572);
sram_add_entry(0, 3, 768, 4, 128'h4030000000000000000c90d419a);
sram_add_entry(0, 3, 772, 4, 128'h4030000000000000000ff7786b6);
sram_add_entry(0, 3, 776, 4, 128'h4030000000000000000694627e0);
sram_add_entry(0, 3, 780, 4, 128'h4030000000000000000509ecf3e);
sram_add_entry(0, 3, 784, 4, 128'h403000000000000000036c22061);
sram_add_entry(0, 3, 788, 4, 128'h40300000000000000006df4f696);
sram_add_entry(0, 3, 792, 4, 128'h403000000000000000036031f0a);
sram_add_entry(0, 3, 796, 4, 128'h40300000000000000000a146f76);
sram_add_entry(0, 3, 800, 4, 128'h4030000000000000000da603da4);
sram_add_entry(0, 3, 804, 4, 128'h40300000000000000001bd1cc16);
sram_add_entry(0, 3, 808, 4, 128'h4030000000000000000b7e843f9);
sram_add_entry(0, 3, 812, 4, 128'h40300000000000000000ba2d6f7);
sram_add_entry(0, 3, 816, 4, 128'h403000000000000000051de637b);
sram_add_entry(0, 3, 820, 4, 128'h4030000000000000000828ec475);
sram_add_entry(0, 3, 824, 4, 128'h4030000000000000000cf441982);
sram_add_entry(0, 3, 828, 4, 128'h40300000000000000006f845ae7);
sram_add_entry(0, 3, 832, 4, 128'h403000000000000000086e14992);
sram_add_entry(0, 3, 836, 4, 128'h4030000000000000000c785a77a);
sram_add_entry(0, 3, 840, 4, 128'h4030000000000000000f41488dc);
sram_add_entry(0, 3, 844, 4, 128'h4030000000000000000dc6d7d76);
sram_add_entry(0, 3, 848, 4, 128'h4030000000000000000b9305c01);
sram_add_entry(0, 3, 852, 4, 128'h40300000000000000001b750d7d);
sram_add_entry(0, 3, 856, 4, 128'h403000000000000000052e6d13c);
sram_add_entry(0, 3, 860, 4, 128'h4030000000000000000c8ae7d5e);
sram_add_entry(0, 3, 864, 4, 128'h4030000000000000000ed2db3be);
sram_add_entry(0, 3, 868, 4, 128'h403000000000000000066f59500);
sram_add_entry(0, 3, 872, 4, 128'h403000000000000000090d448e9);
sram_add_entry(0, 3, 876, 4, 128'h4030000000000000000b51cbc38);
sram_add_entry(0, 3, 880, 4, 128'h403000000000000000047180bae);
sram_add_entry(0, 3, 884, 4, 128'h4030000000000000000e1ffb22b);
sram_add_entry(0, 3, 888, 4, 128'h4030000000000000000eb5391a7);
sram_add_entry(0, 3, 892, 4, 128'h40300000000000000001c9a36cd);
sram_add_entry(0, 3, 896, 4, 128'h40300000000000000009d48a1ec);
sram_add_entry(0, 3, 900, 4, 128'h40300000000000000005163f4bb);
sram_add_entry(0, 3, 904, 4, 128'h403000000000000000063169cd6);
sram_add_entry(0, 3, 908, 4, 128'h4030000000000000000afa075ec);
sram_add_entry(0, 3, 912, 4, 128'h4030000000000000000100c2296);
sram_add_entry(0, 3, 916, 4, 128'h4030000000000000000ee45cc7a);
sram_add_entry(0, 3, 920, 4, 128'h40300000000000000006f92ad29);
sram_add_entry(0, 3, 924, 4, 128'h403000000000000000029b9588d);
sram_add_entry(0, 3, 928, 4, 128'h4030000000000000000618563e7);
sram_add_entry(0, 3, 932, 4, 128'h4030000000000000000a58cb19c);
sram_add_entry(0, 3, 936, 4, 128'h40300000000000000001a5533c0);
sram_add_entry(0, 3, 940, 4, 128'h40300000000000000009afdd7cc);
sram_add_entry(0, 3, 944, 4, 128'h4030000000000000000fb3a8fdc);
sram_add_entry(0, 3, 948, 4, 128'h40300000000000000007739a57a);
sram_add_entry(0, 3, 952, 4, 128'h4030000000000000000bc3079c2);
sram_add_entry(0, 3, 956, 4, 128'h4030000000000000000566dbe9d);
sram_add_entry(0, 3, 960, 4, 128'h4030000000000000000a5b90f20);
sram_add_entry(0, 3, 964, 4, 128'h403000000000000000017bbd94a);
sram_add_entry(0, 3, 968, 4, 128'h4030000000000000000d3cf3d16);
sram_add_entry(0, 3, 972, 4, 128'h40300000000000000004beeacd4);
sram_add_entry(0, 3, 976, 4, 128'h4030000000000000000137474a7);
sram_add_entry(0, 3, 980, 4, 128'h4030000000000000000ec022a40);
sram_add_entry(0, 3, 984, 4, 128'h4030000000000000000a25046c1);
sram_add_entry(0, 3, 988, 4, 128'h40300000000000000007035529d);
sram_add_entry(0, 3, 992, 4, 128'h40300000000000000001cadbeb4);
sram_add_entry(0, 3, 996, 4, 128'h40300000000000000008400df43);
sram_add_entry(0, 3, 1000, 4, 128'h4030000000000000000e6b8086f);
sram_add_entry(0, 3, 1004, 4, 128'h403000000000000000087384f57);
sram_add_entry(0, 3, 1008, 4, 128'h40300000000000000008d078eb8);
sram_add_entry(0, 3, 1012, 4, 128'h4030000000000000000126db093);
sram_add_entry(0, 3, 1016, 4, 128'h4030000000000000000bf6cb612);
sram_add_entry(0, 3, 1020, 4, 128'h4030000000000000000695c7a60);
sram_add_entry(0, 3, 1024, 4, 128'h40300000000000000006c8e6262);
sram_add_entry(0, 3, 1028, 4, 128'h40300000000000000009a4b4a8a);
sram_add_entry(0, 3, 1032, 4, 128'h40300000000000000009dfaf7d0);
sram_add_entry(0, 3, 1036, 4, 128'h403000000000000000022388795);
sram_add_entry(0, 3, 1040, 4, 128'h40300000000000000000706887e);
sram_add_entry(0, 3, 1044, 4, 128'h403000000000000000050674a03);
sram_add_entry(0, 3, 1048, 4, 128'h4030000000000000000c0303373);
sram_add_entry(0, 3, 1052, 4, 128'h4030000000000000000613a337b);
sram_add_entry(0, 3, 1056, 4, 128'h4030000000000000000f56e398f);
sram_add_entry(0, 3, 1060, 4, 128'h403000000000000000076190ad6);
sram_add_entry(0, 3, 1064, 4, 128'h40300000000000000001a074b4d);
sram_add_entry(0, 3, 1068, 4, 128'h4030000000000000000b9d382dd);
sram_add_entry(0, 3, 1072, 4, 128'h403000000000000000049627c77);
sram_add_entry(0, 3, 1076, 4, 128'h40300000000000000001af7fc78);
sram_add_entry(0, 3, 1080, 4, 128'h40300000000000000004c5b58c2);
sram_add_entry(0, 3, 1084, 4, 128'h4030000000000000000f7b90362);
sram_add_entry(0, 3, 1088, 4, 128'h403000000000000000064c19c57);
sram_add_entry(0, 3, 1092, 4, 128'h40300000000000000004ced0ec5);
sram_add_entry(0, 3, 1096, 4, 128'h403000000000000000063da1ff4);
sram_add_entry(0, 3, 1100, 4, 128'h4030000000000000000d2bdc987);
sram_add_entry(0, 3, 1104, 4, 128'h403000000000000000092fa7936);
sram_add_entry(0, 3, 1108, 4, 128'h4030000000000000000f1e9bbdc);
sram_add_entry(0, 3, 1112, 4, 128'h4030000000000000000eb9f570f);
sram_add_entry(0, 3, 1116, 4, 128'h40300000000000000005675f48e);
sram_add_entry(0, 3, 1120, 4, 128'h40300000000000000000e73169c);
sram_add_entry(0, 3, 1124, 4, 128'h403000000000000000012604535);
sram_add_entry(0, 3, 1128, 4, 128'h4030000000000000000f8e3f27b);
sram_add_entry(0, 3, 1132, 4, 128'h4030000000000000000876c9502);
sram_add_entry(0, 3, 1136, 4, 128'h403000000000000000038ecaf18);
sram_add_entry(0, 3, 1140, 4, 128'h403000000000000000010bb22bf);
sram_add_entry(0, 3, 1144, 4, 128'h4030000000000000000f4bef27c);
sram_add_entry(0, 3, 1148, 4, 128'h40300000000000000004cc5a1f3);
sram_add_entry(0, 3, 1152, 4, 128'h4030000000000000000fb03f116);
sram_add_entry(0, 3, 1156, 4, 128'h4030000000000000000001c1d63);
sram_add_entry(0, 3, 1160, 4, 128'h4030000000000000000634ba600);
sram_add_entry(0, 3, 1164, 4, 128'h4030000000000000000b6bfd1ef);
sram_add_entry(0, 3, 1168, 4, 128'h403000000000000000031a5e63f);
sram_add_entry(0, 3, 1172, 4, 128'h4030000000000000000748ba60c);
sram_add_entry(0, 3, 1176, 4, 128'h4030000000000000000642e6f5e);
sram_add_entry(0, 3, 1180, 4, 128'h403000000000000000046f2c3d3);
sram_add_entry(0, 3, 1184, 4, 128'h403000000000000000002636104);
sram_add_entry(0, 3, 1188, 4, 128'h40300000000000000001ebfe132);
sram_add_entry(0, 3, 1192, 4, 128'h40300000000000000002b75c41c);
sram_add_entry(0, 3, 1196, 4, 128'h403000000000000000033c7ddf3);
sram_add_entry(0, 3, 1200, 4, 128'h40300000000000000009d1dd7c9);
sram_add_entry(0, 3, 1204, 4, 128'h403000000000000000056c445e5);
sram_add_entry(0, 3, 1208, 4, 128'h40300000000000000000582da58);
sram_add_entry(0, 3, 1212, 4, 128'h403000000000000000053ea3aa0);
sram_add_entry(0, 3, 1216, 4, 128'h40300000000000000006528ce42);
sram_add_entry(0, 3, 1220, 4, 128'h4030000000000000000a662e2fd);
sram_add_entry(0, 3, 1224, 4, 128'h403000000000000000052fcf82a);
sram_add_entry(0, 3, 1228, 4, 128'h4030000000000000000a36b6724);
sram_add_entry(0, 3, 1232, 4, 128'h403000000000000000057277a34);
sram_add_entry(0, 3, 1236, 4, 128'h40300000000000000008e243f26);
sram_add_entry(0, 3, 1240, 4, 128'h40300000000000000003f9a74c6);
sram_add_entry(0, 3, 1244, 4, 128'h403000000000000000086ae1fea);
sram_add_entry(0, 3, 1248, 4, 128'h403000000000000000009030da8);
sram_add_entry(0, 3, 1252, 4, 128'h4030000000000000000ad1f99b7);
sram_add_entry(0, 3, 1256, 4, 128'h40300000000000000008909580a);
sram_add_entry(0, 3, 1260, 4, 128'h40300000000000000002ec02701);
sram_add_entry(0, 3, 1264, 4, 128'h4030000000000000000397c1787);
sram_add_entry(0, 3, 1268, 4, 128'h403000000000000000018384914);
sram_add_entry(0, 3, 1272, 4, 128'h403000000000000000070844238);
sram_add_entry(0, 3, 1276, 4, 128'h403000000000000000078d836a6);
sram_add_entry(0, 3, 1280, 4, 128'h403000000000000000062a813b2);
sram_add_entry(0, 3, 1284, 4, 128'h4030000000000000000a8218af8);
sram_add_entry(0, 3, 1288, 4, 128'h40300000000000000003fffc90d);
sram_add_entry(0, 3, 1292, 4, 128'h40300000000000000000471270f);
sram_add_entry(0, 3, 1296, 4, 128'h4030000000000000000870c7d6b);
sram_add_entry(0, 3, 1300, 4, 128'h4030000000000000000b1cbd425);
sram_add_entry(0, 3, 1304, 4, 128'h403000000000000000001ca45b7);
sram_add_entry(0, 3, 1308, 4, 128'h4030000000000000000f9b10ce0);
sram_add_entry(0, 3, 1312, 4, 128'h40300000000000000005bc3d7cc);
sram_add_entry(0, 3, 1316, 4, 128'h403000000000000000078b9b3f0);
sram_add_entry(0, 3, 1320, 4, 128'h4030000000000000000d4aa27c8);
sram_add_entry(0, 3, 1324, 4, 128'h40300000000000000005f341aa9);
sram_add_entry(0, 3, 1328, 4, 128'h4030000000000000000ba354357);
sram_add_entry(0, 3, 1332, 4, 128'h403000000000000000088c143b0);
sram_add_entry(0, 3, 1336, 4, 128'h403000000000000000048d9a0b4);
sram_add_entry(0, 3, 1340, 4, 128'h4030000000000000000ab4daf75);
sram_add_entry(0, 3, 1344, 4, 128'h4030000000000000000d975a916);
sram_add_entry(0, 3, 1348, 4, 128'h4030000000000000000e845c902);
sram_add_entry(0, 3, 1352, 4, 128'h4030000000000000000878c2f86);
sram_add_entry(0, 3, 1356, 4, 128'h4030000000000000000ba02f376);
sram_add_entry(0, 3, 1360, 4, 128'h4030000000000000000fe0f25ec);
sram_add_entry(0, 3, 1364, 4, 128'h4030000000000000000bcce8db5);
sram_add_entry(0, 3, 1368, 4, 128'h4030000000000000000c3cb15c5);
sram_add_entry(0, 3, 1372, 4, 128'h403000000000000000032042660);
sram_add_entry(0, 3, 1376, 4, 128'h4030000000000000000713fad01);
sram_add_entry(0, 3, 1380, 4, 128'h40300000000000000001e45babb);
sram_add_entry(0, 3, 1384, 4, 128'h4030000000000000000537ea7b5);
sram_add_entry(0, 3, 1388, 4, 128'h40300000000000000002451b99d);
sram_add_entry(0, 3, 1392, 4, 128'h40300000000000000008c16bba1);
sram_add_entry(0, 3, 1396, 4, 128'h4030000000000000000a6d92913);
sram_add_entry(0, 3, 1400, 4, 128'h4030000000000000000c44e2eee);
sram_add_entry(0, 3, 1404, 4, 128'h40300000000000000009f76d085);
sram_add_entry(0, 3, 1408, 4, 128'h40300000000000000000774bd3b);
sram_add_entry(0, 3, 1412, 4, 128'h4030000000000000000b8c9750b);
sram_add_entry(0, 3, 1416, 4, 128'h40300000000000000003b9ced0c);
sram_add_entry(0, 3, 1420, 4, 128'h4030000000000000000e822c48d);
sram_add_entry(0, 3, 1424, 4, 128'h4030000000000000000605c12f0);
sram_add_entry(0, 3, 1428, 4, 128'h4030000000000000000d1c12819);
sram_add_entry(0, 3, 1432, 4, 128'h403000000000000000048d1d320);
sram_add_entry(0, 3, 1436, 4, 128'h40300000000000000003b2aa084);
sram_add_entry(0, 3, 1440, 4, 128'h403000000000000000016bb4af9);
sram_add_entry(0, 3, 1444, 4, 128'h4030000000000000000fab919eb);
sram_add_entry(0, 3, 1448, 4, 128'h403000000000000000009632817);
sram_add_entry(0, 3, 1452, 4, 128'h40300000000000000002a14c3c5);
sram_add_entry(0, 3, 1456, 4, 128'h4030000000000000000088430aa);
sram_add_entry(0, 3, 1460, 4, 128'h40300000000000000004b138290);
sram_add_entry(0, 3, 1464, 4, 128'h4030000000000000000a4328192);
sram_add_entry(0, 3, 1468, 4, 128'h4030000000000000000af74e5f0);
sram_add_entry(0, 3, 1472, 4, 128'h4030000000000000000adcbcea6);
sram_add_entry(0, 3, 1476, 4, 128'h403000000000000000095e27aa3);
sram_add_entry(0, 3, 1480, 4, 128'h40300000000000000002f201bf5);
sram_add_entry(0, 3, 1484, 4, 128'h4030000000000000000a17dce45);
sram_add_entry(0, 3, 1488, 4, 128'h40300000000000000009267213c);
sram_add_entry(0, 3, 1492, 4, 128'h40300000000000000002307fd2f);
sram_add_entry(0, 3, 1496, 4, 128'h4030000000000000000f7c0c8ec);
sram_add_entry(0, 3, 1500, 4, 128'h4030000000000000000c01c6536);
sram_add_entry(0, 3, 1504, 4, 128'h40300000000000000005821ab3b);
sram_add_entry(0, 3, 1508, 4, 128'h4030000000000000000393a4f1e);
sram_add_entry(0, 3, 1512, 4, 128'h40300000000000000004ccacbaa);
sram_add_entry(0, 3, 1516, 4, 128'h40300000000000000000bb0cce2);
sram_add_entry(0, 3, 1520, 4, 128'h40300000000000000004a3557dc);
sram_add_entry(0, 3, 1524, 4, 128'h4030000000000000000a7f5f126);
sram_add_entry(0, 3, 1528, 4, 128'h4030000000000000000ecbf5817);
sram_add_entry(0, 3, 1532, 4, 128'h40300000000000000004fcce4ae);
sram_add_entry(0, 3, 1536, 4, 128'h403000000000000000049ca82c1);
sram_add_entry(0, 3, 1540, 4, 128'h4030000000000000000c256a85f);
sram_add_entry(0, 3, 1544, 4, 128'h4030000000000000000d0e74b83);
sram_add_entry(0, 3, 1548, 4, 128'h4030000000000000000f790724d);
sram_add_entry(0, 3, 1552, 4, 128'h4030000000000000000aa4fdd5a);
sram_add_entry(0, 3, 1556, 4, 128'h40300000000000000009302e606);
sram_add_entry(0, 3, 1560, 4, 128'h4030000000000000000774c0a95);
sram_add_entry(0, 3, 1564, 4, 128'h4030000000000000000fe7ba7a6);
sram_add_entry(0, 3, 1568, 4, 128'h4030000000000000000763c92c9);
sram_add_entry(0, 3, 1572, 4, 128'h4030000000000000000161007b1);
sram_add_entry(0, 3, 1576, 4, 128'h40300000000000000002a09f69b);
sram_add_entry(0, 3, 1580, 4, 128'h403000000000000000008f0631a);
sram_add_entry(0, 3, 1584, 4, 128'h40300000000000000006e5a5a64);
sram_add_entry(0, 3, 1588, 4, 128'h4030000000000000000e4f1fdf8);
sram_add_entry(0, 3, 1592, 4, 128'h403000000000000000082ee13b8);
sram_add_entry(0, 3, 1596, 4, 128'h40300000000000000003ebac666);
sram_add_entry(0, 3, 1600, 4, 128'h4030000000000000000c30bb880);
sram_add_entry(0, 3, 1604, 4, 128'h40300000000000000007bd0807a);
sram_add_entry(0, 3, 1608, 4, 128'h403000000000000000069c9a36a);
sram_add_entry(0, 3, 1612, 4, 128'h40300000000000000006dfa7ea1);
sram_add_entry(0, 3, 1616, 4, 128'h4030000000000000000465e2174);
sram_add_entry(0, 3, 1620, 4, 128'h4030000000000000000d690c48f);
sram_add_entry(0, 3, 1624, 4, 128'h40300000000000000004dfb8bb3);
sram_add_entry(0, 3, 1628, 4, 128'h4030000000000000000fcfb8a1d);
sram_add_entry(0, 3, 1632, 4, 128'h40300000000000000001e97dfa7);
sram_add_entry(0, 3, 1636, 4, 128'h4030000000000000000fb45ee29);
sram_add_entry(0, 3, 1640, 4, 128'h40300000000000000002e75bd78);
sram_add_entry(0, 3, 1644, 4, 128'h403000000000000000022c82a03);
sram_add_entry(0, 3, 1648, 4, 128'h4030000000000000000b5e57ae6);
sram_add_entry(0, 3, 1652, 4, 128'h40300000000000000006d61818d);
sram_add_entry(0, 3, 1656, 4, 128'h403000000000000000089bd817f);
sram_add_entry(0, 3, 1660, 4, 128'h403000000000000000039a3e363);
sram_add_entry(0, 3, 1664, 4, 128'h4030000000000000000f1d02dcb);
sram_add_entry(0, 3, 1668, 4, 128'h4030000000000000000e7cab4e5);
sram_add_entry(0, 3, 1672, 4, 128'h403000000000000000093c91bc5);
sram_add_entry(0, 3, 1676, 4, 128'h40300000000000000007e18e057);
sram_add_entry(0, 3, 1680, 4, 128'h4030000000000000000a32ff2f6);
sram_add_entry(0, 3, 1684, 4, 128'h4030000000000000000176b62ce);
sram_add_entry(0, 3, 1688, 4, 128'h403000000000000000031482dc2);
sram_add_entry(0, 3, 1692, 4, 128'h40300000000000000005dd0192c);
sram_add_entry(0, 3, 1696, 4, 128'h40300000000000000009c37fed2);
sram_add_entry(0, 3, 1700, 4, 128'h40300000000000000004172ae7a);
sram_add_entry(0, 3, 1704, 4, 128'h40300000000000000007a4b700b);
sram_add_entry(0, 3, 1708, 4, 128'h40300000000000000005b6bae30);
sram_add_entry(0, 3, 1712, 4, 128'h4030000000000000000c829489d);
sram_add_entry(0, 3, 1716, 4, 128'h40300000000000000001fe9c4aa);
sram_add_entry(0, 3, 1720, 4, 128'h4030000000000000000455925b1);
sram_add_entry(0, 3, 1724, 4, 128'h4030000000000000000eec3172f);
sram_add_entry(0, 3, 1728, 4, 128'h4030000000000000000be5b95ba);
sram_add_entry(0, 3, 1732, 4, 128'h4030000000000000000f7c5318d);
sram_add_entry(0, 3, 1736, 4, 128'h403000000000000000032b3ab3d);
sram_add_entry(0, 3, 1740, 4, 128'h4030000000000000000f03288ba);
sram_add_entry(0, 3, 1744, 4, 128'h403000000000000000054d26dab);
sram_add_entry(0, 3, 1748, 4, 128'h40300000000000000003b35ba0b);
sram_add_entry(0, 3, 1752, 4, 128'h40300000000000000004725d7df);
sram_add_entry(0, 3, 1756, 4, 128'h403000000000000000082bd2740);
sram_add_entry(0, 3, 1760, 4, 128'h40300000000000000004ab16fe6);
sram_add_entry(0, 3, 1764, 4, 128'h4030000000000000000b8828761);
sram_add_entry(0, 3, 1768, 4, 128'h4030000000000000000d7fed41e);
sram_add_entry(0, 3, 1772, 4, 128'h4030000000000000000927e89c8);
sram_add_entry(0, 3, 1776, 4, 128'h403000000000000000069ce648c);
sram_add_entry(0, 3, 1780, 4, 128'h4030000000000000000a98af6be);
sram_add_entry(0, 3, 1784, 4, 128'h4030000000000000000830c2297);
sram_add_entry(0, 3, 1788, 4, 128'h40300000000000000008a7c096a);
sram_add_entry(0, 3, 1792, 4, 128'h403000000000000000087b80521);
sram_add_entry(0, 3, 1796, 4, 128'h40300000000000000007b3a4eaa);
sram_add_entry(0, 3, 1800, 4, 128'h4030000000000000000be3050db);
sram_add_entry(0, 3, 1804, 4, 128'h4030000000000000000dc28e522);
sram_add_entry(0, 3, 1808, 4, 128'h403000000000000000036b04f1c);
sram_add_entry(0, 3, 1812, 4, 128'h4030000000000000000403a7c3e);
sram_add_entry(0, 3, 1816, 4, 128'h403000000000000000003955090);
sram_add_entry(0, 3, 1820, 4, 128'h403000000000000000009b0e15b);
sram_add_entry(0, 3, 1824, 4, 128'h40300000000000000009d7eb941);
sram_add_entry(0, 3, 1828, 4, 128'h403000000000000000092cc7b97);
sram_add_entry(0, 3, 1832, 4, 128'h4030000000000000000526e091b);
sram_add_entry(0, 3, 1836, 4, 128'h40300000000000000003f5d769e);
sram_add_entry(0, 3, 1840, 4, 128'h4030000000000000000150c92e2);
sram_add_entry(0, 3, 1844, 4, 128'h4030000000000000000e834138a);
sram_add_entry(0, 3, 1848, 4, 128'h4030000000000000000c34ca9d1);
sram_add_entry(0, 3, 1852, 4, 128'h4030000000000000000b3572efe);
sram_add_entry(0, 3, 1856, 4, 128'h4030000000000000000c6f229f9);
sram_add_entry(0, 3, 1860, 4, 128'h4030000000000000000e5cbabe9);
sram_add_entry(0, 3, 1864, 4, 128'h4030000000000000000864f25f7);
sram_add_entry(0, 3, 1868, 4, 128'h403000000000000000067c4066d);
sram_add_entry(0, 3, 1872, 4, 128'h40300000000000000009de1cb00);
sram_add_entry(0, 3, 1876, 4, 128'h403000000000000000034248c05);
sram_add_entry(0, 3, 1880, 4, 128'h4030000000000000000c58b25e4);
sram_add_entry(0, 3, 1884, 4, 128'h4030000000000000000b3f968f6);
sram_add_entry(0, 3, 1888, 4, 128'h40300000000000000008948dfa0);
sram_add_entry(0, 3, 1892, 4, 128'h40300000000000000006186b4d5);
sram_add_entry(0, 3, 1896, 4, 128'h4030000000000000000e5423ca6);
sram_add_entry(0, 3, 1900, 4, 128'h4030000000000000000fb755c87);
sram_add_entry(0, 3, 1904, 4, 128'h4030000000000000000a2792929);
sram_add_entry(0, 3, 1908, 4, 128'h4030000000000000000d4bca2bb);
sram_add_entry(0, 3, 1912, 4, 128'h40300000000000000003c15896e);
sram_add_entry(0, 3, 1916, 4, 128'h403000000000000000088e915d3);
sram_add_entry(0, 3, 1920, 4, 128'h403000000000000000062db80d6);
sram_add_entry(0, 3, 1924, 4, 128'h40300000000000000004c481bbc);
sram_add_entry(0, 3, 1928, 4, 128'h403000000000000000009dbbbd6);
sram_add_entry(0, 3, 1932, 4, 128'h4030000000000000000fcce66eb);
sram_add_entry(0, 3, 1936, 4, 128'h40300000000000000006830b811);
sram_add_entry(0, 3, 1940, 4, 128'h40300000000000000004379b461);
sram_add_entry(0, 3, 1944, 4, 128'h403000000000000000068938af3);
sram_add_entry(0, 3, 1948, 4, 128'h40300000000000000007ff6250d);
sram_add_entry(0, 3, 1952, 4, 128'h4030000000000000000d0b2e426);
sram_add_entry(0, 3, 1956, 4, 128'h4030000000000000000e0769eb3);
sram_add_entry(0, 3, 1960, 4, 128'h4030000000000000000ebca488e);
sram_add_entry(0, 3, 1964, 4, 128'h4030000000000000000a7d59609);
sram_add_entry(0, 3, 1968, 4, 128'h4030000000000000000861d983b);
sram_add_entry(0, 3, 1972, 4, 128'h403000000000000000013c0f8ae);
sram_add_entry(0, 3, 1976, 4, 128'h40300000000000000009aac6fda);
sram_add_entry(0, 3, 1980, 4, 128'h403000000000000000043d9df1c);
sram_add_entry(0, 3, 1984, 4, 128'h4030000000000000000e9a06c24);
sram_add_entry(0, 3, 1988, 4, 128'h4030000000000000000ac0241b2);
sram_add_entry(0, 3, 1992, 4, 128'h40300000000000000007612253b);
sram_add_entry(0, 3, 1996, 4, 128'h4030000000000000000ed8abb5c);
sram_add_entry(0, 3, 2000, 4, 128'h40300000000000000006f9d5e51);
sram_add_entry(0, 3, 2004, 4, 128'h403000000000000000016ac4efe);
sram_add_entry(0, 3, 2008, 4, 128'h4030000000000000000c3ab0255);
sram_add_entry(0, 3, 2012, 4, 128'h4030000000000000000c4f30409);
sram_add_entry(0, 3, 2016, 4, 128'h403000000000000000039a47d32);
sram_add_entry(0, 3, 2020, 4, 128'h4030000000000000000935c5f96);
sram_add_entry(0, 3, 2024, 4, 128'h403000000000000000046b4c54a);
sram_add_entry(0, 3, 2028, 4, 128'h403000000000000000094b72783);
sram_add_entry(0, 3, 2032, 4, 128'h4030000000000000000b1299113);
sram_add_entry(0, 3, 2036, 4, 128'h40300000000000000008bed837b);
sram_add_entry(0, 3, 2040, 4, 128'h40300000000000000004420d131);
sram_add_entry(0, 3, 2044, 4, 128'h403000000000000000053eb678a);
sram_add_entry(0, 3, 2048, 4, 128'h4030000000000000000bae75dd5);
sram_add_entry(0, 3, 2052, 4, 128'h403000000000000000018f29af4);
sram_add_entry(0, 3, 2056, 4, 128'h403000000000000000034bf20e6);
sram_add_entry(0, 3, 2060, 4, 128'h4030000000000000000d7e1bf9e);
sram_add_entry(0, 3, 2064, 4, 128'h4030000000000000000c653b4a2);
sram_add_entry(0, 3, 2068, 4, 128'h40300000000000000001017a7ee);
sram_add_entry(0, 3, 2072, 4, 128'h40300000000000000007f128a80);
sram_add_entry(0, 3, 2076, 4, 128'h40300000000000000007c5925b4);
sram_add_entry(0, 3, 2080, 4, 128'h40300000000000000004538f048);
sram_add_entry(0, 3, 2084, 4, 128'h4030000000000000000a93c8da7);
sram_add_entry(0, 3, 2088, 4, 128'h4030000000000000000ac4a08d6);
sram_add_entry(0, 3, 2092, 4, 128'h40300000000000000009a0f4cf3);
sram_add_entry(0, 3, 2096, 4, 128'h4030000000000000000f277f763);
sram_add_entry(0, 3, 2100, 4, 128'h40300000000000000008582cf49);
sram_add_entry(0, 3, 2104, 4, 128'h403000000000000000093c3f421);
sram_add_entry(0, 3, 2108, 4, 128'h4030000000000000000918c2423);
sram_add_entry(0, 3, 2112, 4, 128'h40300000000000000009a777ce4);
sram_add_entry(0, 3, 2116, 4, 128'h403000000000000000036dfd172);
sram_add_entry(0, 3, 2120, 4, 128'h4030000000000000000d5556de3);
sram_add_entry(0, 3, 2124, 4, 128'h4030000000000000000ce40b138);
sram_add_entry(0, 3, 2128, 4, 128'h40300000000000000004aeecfc5);
sram_add_entry(0, 3, 2132, 4, 128'h403000000000000000003b5012c);
sram_add_entry(0, 3, 2136, 4, 128'h4030000000000000000a397b379);
sram_add_entry(0, 3, 2140, 4, 128'h4030000000000000000c8efbd35);
sram_add_entry(0, 3, 2144, 4, 128'h4030000000000000000197ecb0c);
sram_add_entry(0, 3, 2148, 4, 128'h40300000000000000003bb510bf);
sram_add_entry(0, 3, 2152, 4, 128'h4030000000000000000c6f6d63e);
sram_add_entry(0, 3, 2156, 4, 128'h4030000000000000000071d6384);
sram_add_entry(0, 3, 2160, 4, 128'h4030000000000000000c552dd1e);
sram_add_entry(0, 3, 2164, 4, 128'h4030000000000000000e643bc17);
sram_add_entry(0, 3, 2168, 4, 128'h403000000000000000043446e4c);
sram_add_entry(0, 3, 2172, 4, 128'h4030000000000000000bcd07cdb);
sram_add_entry(0, 3, 2176, 4, 128'h40300000000000000007cf14608);
sram_add_entry(0, 3, 2180, 4, 128'h4030000000000000000aff02839);
sram_add_entry(0, 3, 2184, 4, 128'h4030000000000000000b6b7b376);
sram_add_entry(0, 3, 2188, 4, 128'h40300000000000000000511eed1);
sram_add_entry(0, 3, 2192, 4, 128'h40300000000000000006485e04d);
sram_add_entry(0, 3, 2196, 4, 128'h4030000000000000000fb48439e);
sram_add_entry(0, 3, 2200, 4, 128'h40300000000000000001fb6623a);
sram_add_entry(0, 3, 2204, 4, 128'h4030000000000000000748d035f);
sram_add_entry(0, 3, 2208, 4, 128'h4030000000000000000f999c215);
sram_add_entry(0, 3, 2212, 4, 128'h403000000000000000036e773ee);
sram_add_entry(0, 3, 2216, 4, 128'h40300000000000000000ccdabd4);
sram_add_entry(0, 3, 2220, 4, 128'h4030000000000000000b9bbdeca);
sram_add_entry(0, 3, 2224, 4, 128'h4030000000000000000ed764ab2);
sram_add_entry(0, 3, 2228, 4, 128'h403000000000000000048bac8d7);
sram_add_entry(0, 3, 2232, 4, 128'h40300000000000000007c5d1f7c);
sram_add_entry(0, 3, 2236, 4, 128'h4030000000000000000b4ce443a);
sram_add_entry(0, 3, 2240, 4, 128'h403000000000000000065f523a7);
sram_add_entry(0, 3, 2244, 4, 128'h40300000000000000007875ba6d);
sram_add_entry(0, 3, 2248, 4, 128'h4030000000000000000c13082b4);
sram_add_entry(0, 3, 2252, 4, 128'h4030000000000000000c606c212);
sram_add_entry(0, 3, 2256, 4, 128'h40300000000000000001e7bb588);
sram_add_entry(0, 3, 2260, 4, 128'h4030000000000000000c05f13a2);
sram_add_entry(0, 3, 2264, 4, 128'h4030000000000000000a10fdd47);
sram_add_entry(0, 3, 2268, 4, 128'h40300000000000000002cd17cd7);
sram_add_entry(0, 3, 2272, 4, 128'h4030000000000000000116e1259);
sram_add_entry(0, 3, 2276, 4, 128'h403000000000000000069fd204c);
sram_add_entry(0, 3, 2280, 4, 128'h403000000000000000012118ecd);
sram_add_entry(0, 3, 2284, 4, 128'h403000000000000000044d49085);
sram_add_entry(0, 3, 2288, 4, 128'h4030000000000000000d7748be2);
sram_add_entry(0, 3, 2292, 4, 128'h403000000000000000062dacdb8);
sram_add_entry(0, 3, 2296, 4, 128'h40300000000000000005d114a9b);
sram_add_entry(0, 3, 2300, 4, 128'h4030000000000000000616bc248);
sram_add_entry(0, 3, 2304, 4, 128'h40300000000000000000b723c38);
sram_add_entry(0, 3, 2308, 4, 128'h4030000000000000000ed1fb3c2);
sram_add_entry(0, 3, 2312, 4, 128'h40300000000000000000f845a6c);
sram_add_entry(0, 3, 2316, 4, 128'h4030000000000000000b66c0f85);
sram_add_entry(0, 3, 2320, 4, 128'h4030000000000000000c7600897);
sram_add_entry(0, 3, 2324, 4, 128'h403000000000000000056100184);
sram_add_entry(0, 3, 2328, 4, 128'h40300000000000000006bcfe5d6);
sram_add_entry(0, 3, 2332, 4, 128'h4030000000000000000cc94b9b7);
sram_add_entry(0, 3, 2336, 4, 128'h403000000000000000029e119ed);
sram_add_entry(0, 3, 2340, 4, 128'h4030000000000000000e11bfdf4);
sram_add_entry(0, 3, 2344, 4, 128'h40300000000000000007acacb1f);
sram_add_entry(0, 3, 2348, 4, 128'h4030000000000000000f4956a20);
sram_add_entry(0, 3, 2352, 4, 128'h4030000000000000000d317a971);
sram_add_entry(0, 3, 2356, 4, 128'h403000000000000000002f31121);
sram_add_entry(0, 3, 2360, 4, 128'h40300000000000000003e589763);
sram_add_entry(0, 3, 2364, 4, 128'h403000000000000000005db4743);
sram_add_entry(0, 3, 2368, 4, 128'h4030000000000000000fc1a80cd);
sram_add_entry(0, 3, 2372, 4, 128'h4030000000000000000651ab564);
sram_add_entry(0, 3, 2376, 4, 128'h403000000000000000008de93c3);
sram_add_entry(0, 3, 2380, 4, 128'h40300000000000000000ff37fd0);
sram_add_entry(0, 3, 2384, 4, 128'h40300000000000000009b657d14);
sram_add_entry(0, 3, 2388, 4, 128'h40300000000000000006309ce86);
sram_add_entry(0, 3, 2392, 4, 128'h403000000000000000073716308);
sram_add_entry(0, 3, 2396, 4, 128'h403000000000000000032c93ff2);
sram_add_entry(0, 3, 2400, 4, 128'h403000000000000000007883f6d);
sram_add_entry(0, 3, 2404, 4, 128'h4030000000000000000ef182c05);
sram_add_entry(0, 3, 2408, 4, 128'h403000000000000000005cf3d0b);
sram_add_entry(0, 3, 2412, 4, 128'h4030000000000000000fa76e3ad);
sram_add_entry(0, 3, 2416, 4, 128'h4030000000000000000cbd8e504);
sram_add_entry(0, 3, 2420, 4, 128'h40300000000000000003318e559);
sram_add_entry(0, 3, 2424, 4, 128'h4030000000000000000d2769959);
sram_add_entry(0, 3, 2428, 4, 128'h403000000000000000054a4165e);
sram_add_entry(0, 3, 2432, 4, 128'h4030000000000000000d19e9f70);
sram_add_entry(0, 3, 2436, 4, 128'h4030000000000000000ed963976);
sram_add_entry(0, 3, 2440, 4, 128'h40300000000000000008c534147);
sram_add_entry(0, 3, 2444, 4, 128'h4030000000000000000d654bf6f);
sram_add_entry(0, 3, 2448, 4, 128'h4030000000000000000e8274dc8);
sram_add_entry(0, 3, 2452, 4, 128'h4030000000000000000153e343f);
sram_add_entry(0, 3, 2456, 4, 128'h403000000000000000076ba647c);
sram_add_entry(0, 3, 2460, 4, 128'h4030000000000000000a78d55ad);
sram_add_entry(0, 3, 2464, 4, 128'h403000000000000000085bef76c);
sram_add_entry(0, 3, 2468, 4, 128'h40300000000000000006b8bdd0e);
sram_add_entry(0, 3, 2472, 4, 128'h40300000000000000003b772627);
sram_add_entry(0, 3, 2476, 4, 128'h40300000000000000009af419a9);
sram_add_entry(0, 3, 2480, 4, 128'h403000000000000000033d61638);
sram_add_entry(0, 3, 2484, 4, 128'h4030000000000000000e0ce4665);
sram_add_entry(0, 3, 2488, 4, 128'h40300000000000000001a783a1f);
sram_add_entry(0, 3, 2492, 4, 128'h40300000000000000000c400047);
sram_add_entry(0, 3, 2496, 4, 128'h4030000000000000000efe82a33);
sram_add_entry(0, 3, 2500, 4, 128'h403000000000000000008fcd729);
sram_add_entry(0, 3, 2504, 4, 128'h4030000000000000000162a2ada);
sram_add_entry(0, 3, 2508, 4, 128'h4030000000000000000a7680901);
sram_add_entry(0, 3, 2512, 4, 128'h4030000000000000000190f7752);
sram_add_entry(0, 3, 2516, 4, 128'h4030000000000000000b6384ac6);
sram_add_entry(0, 3, 2520, 4, 128'h4030000000000000000bbfe5b83);
sram_add_entry(0, 3, 2524, 4, 128'h4030000000000000000cf156c1b);
sram_add_entry(0, 3, 2528, 4, 128'h4030000000000000000da14e4b9);
sram_add_entry(0, 3, 2532, 4, 128'h4030000000000000000f4016e61);
sram_add_entry(0, 3, 2536, 4, 128'h403000000000000000042f4085d);
sram_add_entry(0, 3, 2540, 4, 128'h40300000000000000005ea8c2bd);
sram_add_entry(0, 3, 2544, 4, 128'h4030000000000000000303a3b57);
sram_add_entry(0, 3, 2548, 4, 128'h4030000000000000000b7a150b1);
sram_add_entry(0, 3, 2552, 4, 128'h4030000000000000000fb614d0b);
sram_add_entry(0, 3, 2556, 4, 128'h4030000000000000000e53edcc3);
sram_add_entry(0, 3, 2560, 4, 128'h40300000000000000005b0d54c3);
sram_add_entry(0, 3, 2564, 4, 128'h4030000000000000000605ad057);
sram_add_entry(0, 3, 2568, 4, 128'h40300000000000000008a72fbfe);
sram_add_entry(0, 3, 2572, 4, 128'h40300000000000000004301aa33);
sram_add_entry(0, 3, 2576, 4, 128'h4030000000000000000a29d6bce);
sram_add_entry(0, 3, 2580, 4, 128'h4030000000000000000c2c68789);
sram_add_entry(0, 3, 2584, 4, 128'h40300000000000000007370ec2b);
sram_add_entry(0, 3, 2588, 4, 128'h40300000000000000006989416b);
sram_add_entry(0, 3, 2592, 4, 128'h40300000000000000006f12824b);
sram_add_entry(0, 3, 2596, 4, 128'h403000000000000000021ef3f54);
sram_add_entry(0, 3, 2600, 4, 128'h4030000000000000000b9cd2cd9);
sram_add_entry(0, 3, 2604, 4, 128'h4030000000000000000c0e42d17);
sram_add_entry(0, 3, 2608, 4, 128'h403000000000000000030752c11);
sram_add_entry(0, 3, 2612, 4, 128'h4030000000000000000f36147de);
sram_add_entry(0, 3, 2616, 4, 128'h4030000000000000000dbc68a37);
sram_add_entry(0, 3, 2620, 4, 128'h403000000000000000077949c5f);
sram_add_entry(0, 3, 2624, 4, 128'h4030000000000000000d4ced086);
sram_add_entry(0, 3, 2628, 4, 128'h4030000000000000000f8b6e64c);
sram_add_entry(0, 3, 2632, 4, 128'h403000000000000000044618892);
sram_add_entry(0, 3, 2636, 4, 128'h4030000000000000000bcb45bad);
sram_add_entry(0, 3, 2640, 4, 128'h4030000000000000000da6ce781);
sram_add_entry(0, 3, 2644, 4, 128'h40300000000000000000d3268b7);
sram_add_entry(0, 3, 2648, 4, 128'h4030000000000000000b45e9e05);
sram_add_entry(0, 3, 2652, 4, 128'h4030000000000000000cb3466e1);
sram_add_entry(0, 3, 2656, 4, 128'h4030000000000000000343705e1);
sram_add_entry(0, 3, 2660, 4, 128'h4030000000000000000f235af9a);
sram_add_entry(0, 3, 2664, 4, 128'h4030000000000000000740ad0a0);
sram_add_entry(0, 3, 2668, 4, 128'h4030000000000000000e7680fcb);
sram_add_entry(0, 3, 2672, 4, 128'h4030000000000000000d1ea0b9b);
sram_add_entry(0, 3, 2676, 4, 128'h40300000000000000004e15f57c);
sram_add_entry(0, 3, 2680, 4, 128'h4030000000000000000c059765f);
sram_add_entry(0, 3, 2684, 4, 128'h40300000000000000009df097da);
sram_add_entry(0, 3, 2688, 4, 128'h4030000000000000000c6549881);
sram_add_entry(0, 3, 2692, 4, 128'h4030000000000000000895b90ac);
sram_add_entry(0, 3, 2696, 4, 128'h403000000000000000041466398);
sram_add_entry(0, 3, 2700, 4, 128'h4030000000000000000c6a8e81e);
sram_add_entry(0, 3, 2704, 4, 128'h403000000000000000093ab9460);
sram_add_entry(0, 3, 2708, 4, 128'h4030000000000000000e90e7140);
sram_add_entry(0, 3, 2712, 4, 128'h4030000000000000000f8fb4acb);
sram_add_entry(0, 3, 2716, 4, 128'h40300000000000000001031b5dd);
sram_add_entry(0, 3, 2720, 4, 128'h4030000000000000000e4dc251b);
sram_add_entry(0, 3, 2724, 4, 128'h403000000000000000053d482fa);
sram_add_entry(0, 3, 2728, 4, 128'h4030000000000000000e0ff78f3);
sram_add_entry(0, 3, 2732, 4, 128'h40300000000000000001af2f077);
sram_add_entry(0, 3, 2736, 4, 128'h40300000000000000007bdb5913);
sram_add_entry(0, 3, 2740, 4, 128'h40300000000000000008f40dddc);
sram_add_entry(0, 3, 2744, 4, 128'h403000000000000000017f3c692);
sram_add_entry(0, 3, 2748, 4, 128'h403000000000000000075db959a);
sram_add_entry(0, 3, 2752, 4, 128'h4030000000000000000755727cf);
sram_add_entry(0, 3, 2756, 4, 128'h4030000000000000000374bbaf3);
sram_add_entry(0, 3, 2760, 4, 128'h40300000000000000008a7eca48);
sram_add_entry(0, 3, 2764, 4, 128'h403000000000000000075d671e7);
sram_add_entry(0, 3, 2768, 4, 128'h4030000000000000000f026b004);
sram_add_entry(0, 3, 2772, 4, 128'h4030000000000000000d482915d);
sram_add_entry(0, 3, 2776, 4, 128'h4030000000000000000ee8ec632);
sram_add_entry(0, 3, 2780, 4, 128'h40300000000000000002a2556b1);
sram_add_entry(0, 3, 2784, 4, 128'h40300000000000000003aa3da2c);
sram_add_entry(0, 3, 2788, 4, 128'h403000000000000000062e599fd);
sram_add_entry(0, 3, 2792, 4, 128'h40300000000000000003ad006a9);
sram_add_entry(0, 3, 2796, 4, 128'h40300000000000000000f129a13);
sram_add_entry(0, 3, 2800, 4, 128'h4030000000000000000bd3eb75c);
sram_add_entry(0, 5, 0, 4, 128'h7ab000000000000000000deadbf);
sram_add_entry(0, 5, 4, 4, 128'h40300000000000000005b391854);
sram_add_entry(0, 5, 8, 4, 128'h40300000000000000003e47f882);
sram_add_entry(0, 5, 12, 4, 128'h40300000000000000005914e02b);
sram_add_entry(0, 5, 16, 4, 128'h40300000000000000004195b117);
sram_add_entry(0, 5, 20, 4, 128'h403000000000000000066a71524);
sram_add_entry(0, 5, 24, 4, 128'h403000000000000000051451b67);
sram_add_entry(0, 5, 28, 4, 128'h403000000000000000021189ffb);
sram_add_entry(0, 5, 32, 4, 128'h4030000000000000000cbc0b312);
sram_add_entry(0, 5, 36, 4, 128'h40300000000000000002d22c053);
sram_add_entry(0, 5, 40, 4, 128'h4030000000000000000b3cdad1c);
sram_add_entry(0, 5, 44, 4, 128'h4030000000000000000f1426fee);
sram_add_entry(0, 5, 48, 4, 128'h403000000000000000058f695e9);
sram_add_entry(0, 5, 52, 4, 128'h40300000000000000008c8a5f2f);
sram_add_entry(0, 5, 56, 4, 128'h4030000000000000000a4687d04);
sram_add_entry(0, 5, 60, 4, 128'h4030000000000000000cda417ee);
sram_add_entry(0, 5, 64, 4, 128'h4030000000000000000cc1a14c9);
sram_add_entry(0, 5, 68, 4, 128'h4030000000000000000da52651a);
sram_add_entry(0, 5, 72, 4, 128'h403000000000000000086df7509);
sram_add_entry(0, 5, 76, 4, 128'h40300000000000000004d81cf6e);
sram_add_entry(0, 5, 80, 4, 128'h4030000000000000000bbe63f40);
sram_add_entry(0, 5, 84, 4, 128'h4030000000000000000a2d47841);
sram_add_entry(0, 5, 88, 4, 128'h403000000000000000024aa1d23);
sram_add_entry(0, 5, 92, 4, 128'h403000000000000000083a28630);
sram_add_entry(0, 5, 96, 4, 128'h40300000000000000000f752362);
sram_add_entry(0, 5, 100, 4, 128'h4030000000000000000cf1da1db);
sram_add_entry(0, 5, 104, 4, 128'h403000000000000000005355e83);
sram_add_entry(0, 5, 108, 4, 128'h4030000000000000000b96a09bb);
sram_add_entry(0, 5, 112, 4, 128'h4030000000000000000c02936d5);
sram_add_entry(0, 5, 116, 4, 128'h40300000000000000005d6d63e1);
sram_add_entry(0, 5, 120, 4, 128'h4030000000000000000fbf7c266);
sram_add_entry(0, 5, 124, 4, 128'h4030000000000000000b357e4e5);
sram_add_entry(0, 5, 128, 4, 128'h40300000000000000009b1fb39b);
sram_add_entry(0, 5, 132, 4, 128'h403000000000000000052fb9bde);
sram_add_entry(0, 5, 136, 4, 128'h4030000000000000000fca1984d);
sram_add_entry(0, 5, 140, 4, 128'h4030000000000000000740649d4);
sram_add_entry(0, 5, 144, 4, 128'h40300000000000000009fe5838f);
sram_add_entry(0, 5, 148, 4, 128'h4030000000000000000d0e352d5);
sram_add_entry(0, 5, 152, 4, 128'h4030000000000000000ec62b4dc);
sram_add_entry(0, 5, 156, 4, 128'h4030000000000000000c36e613b);
sram_add_entry(0, 5, 160, 4, 128'h4030000000000000000005479fe);
sram_add_entry(0, 5, 164, 4, 128'h4030000000000000000dbd26ba9);
sram_add_entry(0, 5, 168, 4, 128'h4030000000000000000d6df9413);
sram_add_entry(0, 5, 172, 4, 128'h4030000000000000000c385e52b);
sram_add_entry(0, 5, 176, 4, 128'h4030000000000000000c476407e);
sram_add_entry(0, 5, 180, 4, 128'h403000000000000000025bb9adf);
sram_add_entry(0, 5, 184, 4, 128'h4030000000000000000afef0d47);
sram_add_entry(0, 5, 188, 4, 128'h40300000000000000001b798fdf);
sram_add_entry(0, 5, 192, 4, 128'h403000000000000000031a3da4a);
sram_add_entry(0, 5, 196, 4, 128'h4030000000000000000c5ed41ab);
sram_add_entry(0, 5, 200, 4, 128'h4030000000000000000ba3cc864);
sram_add_entry(0, 5, 204, 4, 128'h403000000000000000032ef62f2);
sram_add_entry(0, 5, 208, 4, 128'h40300000000000000006c4301a5);
sram_add_entry(0, 5, 212, 4, 128'h4030000000000000000235a7415);
sram_add_entry(0, 5, 216, 4, 128'h4030000000000000000e83475e2);
sram_add_entry(0, 5, 220, 4, 128'h40300000000000000005efe85e6);
sram_add_entry(0, 5, 224, 4, 128'h4030000000000000000bb4b49f8);
sram_add_entry(0, 5, 228, 4, 128'h4030000000000000000df9df74d);
sram_add_entry(0, 5, 232, 4, 128'h40300000000000000006633fdf5);
sram_add_entry(0, 5, 236, 4, 128'h4030000000000000000271dda58);
sram_add_entry(0, 5, 240, 4, 128'h40300000000000000003b9537e2);
sram_add_entry(0, 5, 244, 4, 128'h4030000000000000000029f59cc);
sram_add_entry(0, 5, 248, 4, 128'h4030000000000000000214f6a30);
sram_add_entry(0, 5, 252, 4, 128'h4030000000000000000301509db);
sram_add_entry(0, 5, 256, 4, 128'h40300000000000000009675af7b);
sram_add_entry(0, 5, 260, 4, 128'h4030000000000000000623a5d56);
sram_add_entry(0, 5, 264, 4, 128'h4030000000000000000b072e20e);
sram_add_entry(0, 5, 268, 4, 128'h4030000000000000000ff1ffbde);
sram_add_entry(0, 5, 272, 4, 128'h4030000000000000000e73e0b0f);
sram_add_entry(0, 5, 276, 4, 128'h4030000000000000000142ef689);
sram_add_entry(0, 5, 280, 4, 128'h4030000000000000000f1aaddea);
sram_add_entry(0, 5, 284, 4, 128'h403000000000000000052626454);
sram_add_entry(0, 5, 288, 4, 128'h4030000000000000000a731740c);
sram_add_entry(0, 5, 292, 4, 128'h403000000000000000091de6f55);
sram_add_entry(0, 5, 296, 4, 128'h40300000000000000003ae6fcaa);
sram_add_entry(0, 5, 300, 4, 128'h40300000000000000006d454300);
sram_add_entry(0, 5, 304, 4, 128'h403000000000000000044403806);
sram_add_entry(0, 5, 308, 4, 128'h403000000000000000090a17056);
sram_add_entry(0, 5, 312, 4, 128'h4030000000000000000d6246cf5);
sram_add_entry(0, 5, 316, 4, 128'h403000000000000000072c15812);
sram_add_entry(0, 5, 320, 4, 128'h40300000000000000009eac0e5d);
sram_add_entry(0, 5, 324, 4, 128'h4030000000000000000a78d57a7);
sram_add_entry(0, 5, 328, 4, 128'h4030000000000000000b5fb3b40);
sram_add_entry(0, 5, 332, 4, 128'h4030000000000000000c6d29d2b);
sram_add_entry(0, 5, 336, 4, 128'h4030000000000000000e2e8b161);
sram_add_entry(0, 5, 340, 4, 128'h4030000000000000000c9794b3d);
sram_add_entry(0, 5, 344, 4, 128'h4030000000000000000662da1a8);
sram_add_entry(0, 5, 348, 4, 128'h40300000000000000006642c62e);
sram_add_entry(0, 5, 352, 4, 128'h4030000000000000000a3b6c0c1);
sram_add_entry(0, 5, 356, 4, 128'h4030000000000000000c24d613d);
sram_add_entry(0, 5, 360, 4, 128'h4030000000000000000910917bf);
sram_add_entry(0, 5, 364, 4, 128'h40300000000000000003155f993);
sram_add_entry(0, 5, 368, 4, 128'h40300000000000000002a6f131a);
sram_add_entry(0, 5, 372, 4, 128'h4030000000000000000e3b4b767);
sram_add_entry(0, 5, 376, 4, 128'h4030000000000000000e0ae5572);
sram_add_entry(0, 5, 380, 4, 128'h4030000000000000000a94d69c6);
sram_add_entry(0, 5, 384, 4, 128'h40300000000000000006195fa59);
sram_add_entry(0, 5, 388, 4, 128'h403000000000000000095f69846);
sram_add_entry(0, 5, 392, 4, 128'h4030000000000000000e827b8be);
sram_add_entry(0, 5, 396, 4, 128'h4030000000000000000b8ac9596);
sram_add_entry(0, 5, 400, 4, 128'h40300000000000000000ddf142e);
sram_add_entry(0, 5, 404, 4, 128'h40300000000000000005314b7fd);
sram_add_entry(0, 5, 408, 4, 128'h40300000000000000007ea588c1);
sram_add_entry(0, 5, 412, 4, 128'h4030000000000000000af21ab63);
sram_add_entry(0, 5, 416, 4, 128'h40300000000000000005eb7a1ad);
sram_add_entry(0, 5, 420, 4, 128'h4030000000000000000dccbcdaa);
sram_add_entry(0, 5, 424, 4, 128'h4030000000000000000626ccf1e);
sram_add_entry(0, 5, 428, 4, 128'h403000000000000000046c8d7ad);
sram_add_entry(0, 5, 432, 4, 128'h4030000000000000000b278cf5a);
sram_add_entry(0, 5, 436, 4, 128'h4030000000000000000e34af42a);
sram_add_entry(0, 5, 440, 4, 128'h4030000000000000000c927dedb);
sram_add_entry(0, 5, 444, 4, 128'h4030000000000000000ee6dd01c);
sram_add_entry(0, 5, 448, 4, 128'h4030000000000000000df79afea);
sram_add_entry(0, 5, 452, 4, 128'h4030000000000000000b711e4ad);
sram_add_entry(0, 5, 456, 4, 128'h4030000000000000000525533c2);
sram_add_entry(0, 5, 460, 4, 128'h4030000000000000000bdc263d3);
sram_add_entry(0, 5, 464, 4, 128'h4030000000000000000592e4945);
sram_add_entry(0, 5, 468, 4, 128'h4030000000000000000e9b90599);
sram_add_entry(0, 5, 472, 4, 128'h4030000000000000000956729f4);
sram_add_entry(0, 5, 476, 4, 128'h4030000000000000000f35f3a5e);
sram_add_entry(0, 5, 480, 4, 128'h40300000000000000007ab0f7bc);
sram_add_entry(0, 5, 484, 4, 128'h4030000000000000000638321a1);
sram_add_entry(0, 5, 488, 4, 128'h403000000000000000028e8ce21);
sram_add_entry(0, 5, 492, 4, 128'h403000000000000000058309313);
sram_add_entry(0, 5, 496, 4, 128'h403000000000000000014bac6b5);
sram_add_entry(0, 5, 500, 4, 128'h4030000000000000000262308ed);
sram_add_entry(0, 5, 504, 4, 128'h403000000000000000082928ac6);
sram_add_entry(0, 5, 508, 4, 128'h403000000000000000001fa962b);
sram_add_entry(0, 5, 512, 4, 128'h40300000000000000004530cf55);
sram_add_entry(0, 5, 516, 4, 128'h4030000000000000000b7031fdc);
sram_add_entry(0, 5, 520, 4, 128'h40300000000000000003f72ee54);
sram_add_entry(0, 5, 524, 4, 128'h40300000000000000004aef92a8);
sram_add_entry(0, 5, 528, 4, 128'h40300000000000000007dfb9e62);
sram_add_entry(0, 5, 532, 4, 128'h4030000000000000000fd4d55c0);
sram_add_entry(0, 5, 536, 4, 128'h4030000000000000000df11a902);
sram_add_entry(0, 5, 540, 4, 128'h4030000000000000000a994cec8);
sram_add_entry(0, 5, 544, 4, 128'h40300000000000000008b112348);
sram_add_entry(0, 5, 548, 4, 128'h4030000000000000000c5b510b9);
sram_add_entry(0, 5, 552, 4, 128'h403000000000000000011d4a9aa);
sram_add_entry(0, 5, 556, 4, 128'h4030000000000000000654037d5);
sram_add_entry(0, 5, 560, 4, 128'h4030000000000000000b69b89dc);
sram_add_entry(0, 5, 564, 4, 128'h4030000000000000000d8ece25f);
sram_add_entry(0, 5, 568, 4, 128'h4030000000000000000ef864456);
sram_add_entry(0, 5, 572, 4, 128'h40300000000000000007b94efcc);
sram_add_entry(0, 5, 576, 4, 128'h40300000000000000005f914f66);
sram_add_entry(0, 5, 580, 4, 128'h403000000000000000030cd16e7);
sram_add_entry(0, 5, 584, 4, 128'h40300000000000000006e43f380);
sram_add_entry(0, 5, 588, 4, 128'h4030000000000000000aa9b6cac);
sram_add_entry(0, 5, 592, 4, 128'h4030000000000000000cf4b728d);
sram_add_entry(0, 5, 596, 4, 128'h403000000000000000076fbb46a);
sram_add_entry(0, 5, 600, 4, 128'h4030000000000000000060d90ae);
sram_add_entry(0, 5, 604, 4, 128'h4030000000000000000cd54a04b);
sram_add_entry(0, 5, 608, 4, 128'h4030000000000000000cfe265ce);
sram_add_entry(0, 5, 612, 4, 128'h4030000000000000000f0077206);
sram_add_entry(0, 5, 616, 4, 128'h40300000000000000003dd0f100);
sram_add_entry(0, 5, 620, 4, 128'h4030000000000000000fe370614);
sram_add_entry(0, 5, 624, 4, 128'h403000000000000000086391376);
sram_add_entry(0, 5, 628, 4, 128'h4030000000000000000241d8645);
sram_add_entry(0, 5, 632, 4, 128'h4030000000000000000e054378d);
sram_add_entry(0, 5, 636, 4, 128'h4030000000000000000584787de);
sram_add_entry(0, 5, 640, 4, 128'h40300000000000000000c1d8a74);
sram_add_entry(0, 5, 644, 4, 128'h40300000000000000008552542f);
sram_add_entry(0, 5, 648, 4, 128'h40300000000000000006c061d4c);
sram_add_entry(0, 5, 652, 4, 128'h403000000000000000082c410f7);
sram_add_entry(0, 5, 656, 4, 128'h40300000000000000001b55f2a5);
sram_add_entry(0, 5, 660, 4, 128'h403000000000000000019821382);
sram_add_entry(0, 5, 664, 4, 128'h4030000000000000000fc383767);
sram_add_entry(0, 5, 668, 4, 128'h4030000000000000000261dc3a4);
sram_add_entry(0, 5, 672, 4, 128'h403000000000000000066ecf2c0);
sram_add_entry(0, 5, 676, 4, 128'h403000000000000000052965345);
sram_add_entry(0, 5, 680, 4, 128'h403000000000000000033c3d5ba);
sram_add_entry(0, 5, 684, 4, 128'h40300000000000000003debd5fc);
sram_add_entry(0, 5, 688, 4, 128'h403000000000000000030b16b83);
sram_add_entry(0, 5, 692, 4, 128'h40300000000000000009c363d21);
sram_add_entry(0, 5, 696, 4, 128'h403000000000000000061a9a8d5);
sram_add_entry(0, 5, 700, 4, 128'h40300000000000000007c6464e6);
sram_add_entry(0, 5, 704, 4, 128'h403000000000000000000122eb0);
sram_add_entry(0, 5, 708, 4, 128'h4030000000000000000564d3063);
sram_add_entry(0, 5, 712, 4, 128'h403000000000000000092ace320);
sram_add_entry(0, 5, 716, 4, 128'h4030000000000000000d45a4476);
sram_add_entry(0, 5, 720, 4, 128'h403000000000000000082700c14);
sram_add_entry(0, 5, 724, 4, 128'h403000000000000000051c1fec6);
sram_add_entry(0, 5, 728, 4, 128'h4030000000000000000be3dfa7b);
sram_add_entry(0, 5, 732, 4, 128'h403000000000000000017e20095);
sram_add_entry(0, 5, 736, 4, 128'h4030000000000000000d182ec77);
sram_add_entry(0, 5, 740, 4, 128'h40300000000000000001917b9b3);
sram_add_entry(0, 5, 744, 4, 128'h403000000000000000069a64bf6);
sram_add_entry(0, 5, 748, 4, 128'h4030000000000000000c48d51a9);
sram_add_entry(0, 5, 752, 4, 128'h40300000000000000005a3898ac);
sram_add_entry(0, 5, 756, 4, 128'h4030000000000000000ab1e93a4);
sram_add_entry(0, 5, 760, 4, 128'h4030000000000000000ff34d4ee);
sram_add_entry(0, 5, 764, 4, 128'h4030000000000000000d7ec1785);
sram_add_entry(0, 5, 768, 4, 128'h4030000000000000000f631838c);
sram_add_entry(0, 5, 772, 4, 128'h403000000000000000070b5c77e);
sram_add_entry(0, 5, 776, 4, 128'h4030000000000000000f75cba4e);
sram_add_entry(0, 5, 780, 4, 128'h4030000000000000000aa1de942);
sram_add_entry(0, 5, 784, 4, 128'h403000000000000000081a5c739);
sram_add_entry(0, 5, 788, 4, 128'h403000000000000000099781523);
sram_add_entry(0, 5, 792, 4, 128'h4030000000000000000728f2c47);
sram_add_entry(0, 5, 796, 4, 128'h4030000000000000000caf6348c);
sram_add_entry(0, 5, 800, 4, 128'h4030000000000000000ea9c6e6a);
sram_add_entry(0, 5, 804, 4, 128'h403000000000000000029f7a8b6);
sram_add_entry(0, 5, 808, 4, 128'h4030000000000000000b2b48afc);
sram_add_entry(0, 5, 812, 4, 128'h4030000000000000000007ce2de);
sram_add_entry(0, 5, 816, 4, 128'h4030000000000000000e9399dcc);
sram_add_entry(0, 5, 820, 4, 128'h403000000000000000042d77ee9);
sram_add_entry(0, 5, 824, 4, 128'h40300000000000000003fbab7ac);
sram_add_entry(0, 5, 828, 4, 128'h4030000000000000000d2447ab1);
sram_add_entry(0, 5, 832, 4, 128'h40300000000000000001153bd56);
sram_add_entry(0, 5, 836, 4, 128'h4030000000000000000903d6fbe);
sram_add_entry(0, 5, 840, 4, 128'h4030000000000000000057510c1);
sram_add_entry(0, 5, 844, 4, 128'h4030000000000000000e6ed5c85);
sram_add_entry(0, 5, 848, 4, 128'h4030000000000000000311ca0be);
sram_add_entry(0, 5, 852, 4, 128'h4030000000000000000f7280a93);
sram_add_entry(0, 5, 856, 4, 128'h40300000000000000002e6b5b5c);
sram_add_entry(0, 5, 860, 4, 128'h403000000000000000046919b60);
sram_add_entry(0, 5, 864, 4, 128'h4030000000000000000c582966e);
sram_add_entry(0, 5, 868, 4, 128'h4030000000000000000994201b4);
sram_add_entry(0, 5, 872, 4, 128'h40300000000000000000aa59313);
sram_add_entry(0, 5, 876, 4, 128'h4030000000000000000bf51da19);
sram_add_entry(0, 5, 880, 4, 128'h403000000000000000018fa858a);
sram_add_entry(0, 5, 884, 4, 128'h40300000000000000009af5b012);
sram_add_entry(0, 5, 888, 4, 128'h4030000000000000000fe2e0794);
sram_add_entry(0, 5, 892, 4, 128'h403000000000000000086f6eff0);
sram_add_entry(0, 5, 896, 4, 128'h40300000000000000006db30707);
sram_add_entry(0, 5, 900, 4, 128'h403000000000000000027042389);
sram_add_entry(0, 5, 904, 4, 128'h40300000000000000000018914c);
sram_add_entry(0, 5, 908, 4, 128'h40300000000000000001fe68bc6);
sram_add_entry(0, 5, 912, 4, 128'h4030000000000000000a4cd25e8);
sram_add_entry(0, 5, 916, 4, 128'h40300000000000000009dd2002e);
sram_add_entry(0, 5, 920, 4, 128'h4030000000000000000fc0a0251);
sram_add_entry(0, 5, 924, 4, 128'h40300000000000000003c00e18b);
sram_add_entry(0, 5, 928, 4, 128'h40300000000000000001805c387);
sram_add_entry(0, 5, 932, 4, 128'h40300000000000000004f21587a);
sram_add_entry(0, 5, 936, 4, 128'h4030000000000000000182f28a4);
sram_add_entry(0, 5, 940, 4, 128'h4030000000000000000d1f512d2);
sram_add_entry(0, 5, 944, 4, 128'h4030000000000000000b807c52d);
sram_add_entry(0, 5, 948, 4, 128'h4030000000000000000e29931ca);
sram_add_entry(0, 5, 952, 4, 128'h4030000000000000000ace9bab6);
sram_add_entry(0, 5, 956, 4, 128'h4030000000000000000f553012f);
sram_add_entry(0, 5, 960, 4, 128'h4030000000000000000e71db873);
sram_add_entry(0, 5, 964, 4, 128'h4030000000000000000fa51e2d7);
sram_add_entry(0, 5, 968, 4, 128'h4030000000000000000a2049980);
sram_add_entry(0, 5, 972, 4, 128'h4030000000000000000dcabc03c);
sram_add_entry(0, 5, 976, 4, 128'h40300000000000000000eaba455);
sram_add_entry(0, 5, 980, 4, 128'h4030000000000000000a03e1c48);
sram_add_entry(0, 5, 984, 4, 128'h4030000000000000000bd9737aa);
sram_add_entry(0, 5, 988, 4, 128'h40300000000000000008d5ce6fa);
sram_add_entry(0, 5, 992, 4, 128'h4030000000000000000a332a6c7);
sram_add_entry(0, 5, 996, 4, 128'h4030000000000000000d2d22924);
sram_add_entry(0, 5, 1000, 4, 128'h4030000000000000000db0b6f34);
sram_add_entry(0, 5, 1004, 4, 128'h4030000000000000000205831d3);
sram_add_entry(0, 5, 1008, 4, 128'h40300000000000000003423f5ae);
sram_add_entry(0, 5, 1012, 4, 128'h4030000000000000000f69a827f);
sram_add_entry(0, 5, 1016, 4, 128'h4030000000000000000d96cf06f);
sram_add_entry(0, 5, 1020, 4, 128'h4030000000000000000ab53b800);
sram_add_entry(0, 5, 1024, 4, 128'h403000000000000000023b65e4f);
sram_add_entry(0, 5, 1028, 4, 128'h403000000000000000093aeabfb);
sram_add_entry(0, 5, 1032, 4, 128'h4030000000000000000d6166a86);
sram_add_entry(0, 5, 1036, 4, 128'h403000000000000000014acd40b);
sram_add_entry(0, 5, 1040, 4, 128'h403000000000000000070c7ab10);
sram_add_entry(0, 5, 1044, 4, 128'h403000000000000000085c0749b);
sram_add_entry(0, 5, 1048, 4, 128'h403000000000000000040e49bc4);
sram_add_entry(0, 5, 1052, 4, 128'h4030000000000000000d33d79e6);
sram_add_entry(0, 5, 1056, 4, 128'h403000000000000000069bcc50f);
sram_add_entry(0, 5, 1060, 4, 128'h4030000000000000000102d9dfb);
sram_add_entry(0, 5, 1064, 4, 128'h4030000000000000000d9113f9f);
sram_add_entry(0, 5, 1068, 4, 128'h403000000000000000047b3eb80);
sram_add_entry(0, 5, 1072, 4, 128'h4030000000000000000eebaf9d5);
sram_add_entry(0, 5, 1076, 4, 128'h4030000000000000000ebf5e752);
sram_add_entry(0, 5, 1080, 4, 128'h4030000000000000000c857f0a1);
sram_add_entry(0, 5, 1084, 4, 128'h403000000000000000079cedbd6);
sram_add_entry(0, 5, 1088, 4, 128'h4030000000000000000719f8337);
sram_add_entry(0, 5, 1092, 4, 128'h40300000000000000004932ef53);
sram_add_entry(0, 5, 1096, 4, 128'h403000000000000000079ea4387);
sram_add_entry(0, 5, 1100, 4, 128'h403000000000000000074a43cf4);
sram_add_entry(0, 5, 1104, 4, 128'h40300000000000000004fae7a9c);
sram_add_entry(0, 5, 1108, 4, 128'h4030000000000000000117ccf94);
sram_add_entry(0, 5, 1112, 4, 128'h40300000000000000002009284c);
sram_add_entry(0, 5, 1116, 4, 128'h4030000000000000000fd97e863);
sram_add_entry(0, 5, 1120, 4, 128'h4030000000000000000b4be0194);
sram_add_entry(0, 5, 1124, 4, 128'h4030000000000000000379a4aab);
sram_add_entry(0, 5, 1128, 4, 128'h403000000000000000019c749de);
sram_add_entry(0, 5, 1132, 4, 128'h4030000000000000000409fb84d);
sram_add_entry(0, 5, 1136, 4, 128'h40300000000000000003f53200b);
sram_add_entry(0, 5, 1140, 4, 128'h4030000000000000000f7160cc5);
sram_add_entry(0, 5, 1144, 4, 128'h4030000000000000000f8145fad);
sram_add_entry(0, 5, 1148, 4, 128'h4030000000000000000d19b7ecd);
sram_add_entry(0, 5, 1152, 4, 128'h40300000000000000000bb9956a);
sram_add_entry(0, 5, 1156, 4, 128'h4030000000000000000bfc2e567);
sram_add_entry(0, 5, 1160, 4, 128'h4030000000000000000efe2da10);
sram_add_entry(0, 5, 1164, 4, 128'h40300000000000000008359e399);
sram_add_entry(0, 5, 1168, 4, 128'h40300000000000000008352ddc5);
sram_add_entry(0, 5, 1172, 4, 128'h40300000000000000009a537628);
sram_add_entry(0, 5, 1176, 4, 128'h4030000000000000000e7259ec5);
sram_add_entry(0, 5, 1180, 4, 128'h4030000000000000000a2aa7d6d);
sram_add_entry(0, 5, 1184, 4, 128'h4030000000000000000562cb1c9);
sram_add_entry(0, 5, 1188, 4, 128'h4030000000000000000f3c4a8d4);
sram_add_entry(0, 5, 1192, 4, 128'h403000000000000000092ab903f);
sram_add_entry(0, 5, 1196, 4, 128'h403000000000000000055f5e147);
sram_add_entry(0, 5, 1200, 4, 128'h40300000000000000007a4d1421);
sram_add_entry(0, 5, 1204, 4, 128'h40300000000000000007295d548);
sram_add_entry(0, 5, 1208, 4, 128'h40300000000000000004e27af39);
sram_add_entry(0, 5, 1212, 4, 128'h40300000000000000003cc0f13c);
sram_add_entry(0, 5, 1216, 4, 128'h403000000000000000080598983);
sram_add_entry(0, 5, 1220, 4, 128'h403000000000000000003879539);
sram_add_entry(0, 5, 1224, 4, 128'h4030000000000000000c189aa13);
sram_add_entry(0, 5, 1228, 4, 128'h4030000000000000000c9a30d74);
sram_add_entry(0, 5, 1232, 4, 128'h4030000000000000000a560670f);
sram_add_entry(0, 5, 1236, 4, 128'h40300000000000000007565e7f0);
sram_add_entry(0, 5, 1240, 4, 128'h4030000000000000000629f25ce);
sram_add_entry(0, 5, 1244, 4, 128'h4030000000000000000055a2a3e);
sram_add_entry(0, 5, 1248, 4, 128'h4030000000000000000b0a85a06);
sram_add_entry(0, 5, 1252, 4, 128'h4030000000000000000eeefdd01);
sram_add_entry(0, 5, 1256, 4, 128'h4030000000000000000227ae3eb);
sram_add_entry(0, 5, 1260, 4, 128'h40300000000000000002bbb2043);
sram_add_entry(0, 5, 1264, 4, 128'h40300000000000000007c6161ba);
sram_add_entry(0, 5, 1268, 4, 128'h403000000000000000066da02b6);
sram_add_entry(0, 5, 1272, 4, 128'h40300000000000000002d6e83ce);
sram_add_entry(0, 5, 1276, 4, 128'h40300000000000000005e0ed5fd);
sram_add_entry(0, 5, 1280, 4, 128'h40300000000000000004e41522e);
sram_add_entry(0, 5, 1284, 4, 128'h4030000000000000000d651b46b);
sram_add_entry(0, 5, 1288, 4, 128'h403000000000000000062d1130b);
sram_add_entry(0, 5, 1292, 4, 128'h4030000000000000000d35fc028);
sram_add_entry(0, 5, 1296, 4, 128'h40300000000000000005f77f850);
sram_add_entry(0, 5, 1300, 4, 128'h4030000000000000000f6d659f8);
sram_add_entry(0, 5, 1304, 4, 128'h403000000000000000055963f23);
sram_add_entry(0, 5, 1308, 4, 128'h40300000000000000000d4b3416);
sram_add_entry(0, 5, 1312, 4, 128'h4030000000000000000115c174c);
sram_add_entry(0, 5, 1316, 4, 128'h4030000000000000000c120820c);
sram_add_entry(0, 5, 1320, 4, 128'h4030000000000000000f26eb020);
sram_add_entry(0, 5, 1324, 4, 128'h403000000000000000013329e53);
sram_add_entry(0, 5, 1328, 4, 128'h40300000000000000005b10314d);
sram_add_entry(0, 5, 1332, 4, 128'h40300000000000000001e060ea5);
sram_add_entry(0, 5, 1336, 4, 128'h4030000000000000000ff71e09f);
sram_add_entry(0, 5, 1340, 4, 128'h40300000000000000001f6052ef);
sram_add_entry(0, 5, 1344, 4, 128'h4030000000000000000e74d7298);
sram_add_entry(0, 5, 1348, 4, 128'h40300000000000000006bc68533);
sram_add_entry(0, 5, 1352, 4, 128'h4030000000000000000ac2f4971);
sram_add_entry(0, 5, 1356, 4, 128'h4030000000000000000e09c405c);
sram_add_entry(0, 5, 1360, 4, 128'h40300000000000000000bbcf571);
sram_add_entry(0, 5, 1364, 4, 128'h40300000000000000009cb2baa9);
sram_add_entry(0, 5, 1368, 4, 128'h4030000000000000000f9c5b3ea);
sram_add_entry(0, 5, 1372, 4, 128'h4030000000000000000f650f3be);
sram_add_entry(0, 5, 1376, 4, 128'h4030000000000000000d22e73ae);
sram_add_entry(0, 5, 1380, 4, 128'h4030000000000000000d96940ac);
sram_add_entry(0, 5, 1384, 4, 128'h403000000000000000070cd97c2);
sram_add_entry(0, 5, 1388, 4, 128'h4030000000000000000313273e5);
sram_add_entry(0, 5, 1392, 4, 128'h4030000000000000000e79d22d3);
sram_add_entry(0, 5, 1396, 4, 128'h40300000000000000004542cf7e);
sram_add_entry(0, 5, 1400, 4, 128'h403000000000000000086391c8b);
sram_add_entry(0, 5, 1404, 4, 128'h40300000000000000003d91212e);
sram_add_entry(0, 5, 1408, 4, 128'h4030000000000000000c9c85bde);
sram_add_entry(0, 5, 1412, 4, 128'h4030000000000000000c7acf9d9);
sram_add_entry(0, 5, 1416, 4, 128'h4030000000000000000ca0ddcf5);
sram_add_entry(0, 5, 1420, 4, 128'h4030000000000000000d10700da);
sram_add_entry(0, 5, 1424, 4, 128'h40300000000000000003d5daf6b);
sram_add_entry(0, 5, 1428, 4, 128'h403000000000000000016276984);
sram_add_entry(0, 5, 1432, 4, 128'h40300000000000000001267258a);
sram_add_entry(0, 5, 1436, 4, 128'h4030000000000000000a7935c99);
sram_add_entry(0, 5, 1440, 4, 128'h403000000000000000040d7269d);
sram_add_entry(0, 5, 1444, 4, 128'h40300000000000000003b7070ca);
sram_add_entry(0, 5, 1448, 4, 128'h4030000000000000000a265004e);
sram_add_entry(0, 5, 1452, 4, 128'h403000000000000000005aa3264);
sram_add_entry(0, 5, 1456, 4, 128'h4030000000000000000fc21ce68);
sram_add_entry(0, 5, 1460, 4, 128'h4030000000000000000ee6756c9);
sram_add_entry(0, 5, 1464, 4, 128'h4030000000000000000250a4770);
sram_add_entry(0, 5, 1468, 4, 128'h4030000000000000000bb4715f1);
sram_add_entry(0, 5, 1472, 4, 128'h4030000000000000000257f8471);
sram_add_entry(0, 5, 1476, 4, 128'h4030000000000000000181e4032);
sram_add_entry(0, 5, 1480, 4, 128'h4030000000000000000eba8beed);
sram_add_entry(0, 5, 1484, 4, 128'h4030000000000000000550cbdfd);
sram_add_entry(0, 5, 1488, 4, 128'h4030000000000000000312fd6e0);
sram_add_entry(0, 5, 1492, 4, 128'h403000000000000000051244eaf);
sram_add_entry(0, 5, 1496, 4, 128'h403000000000000000033bdf527);
sram_add_entry(0, 5, 1500, 4, 128'h4030000000000000000d14622c5);
sram_add_entry(0, 5, 1504, 4, 128'h4030000000000000000dc47ec5f);
sram_add_entry(0, 5, 1508, 4, 128'h403000000000000000059ac3723);
sram_add_entry(0, 5, 1512, 4, 128'h4030000000000000000c1e60747);
sram_add_entry(0, 5, 1516, 4, 128'h4030000000000000000f7a199f9);
sram_add_entry(0, 5, 1520, 4, 128'h40300000000000000005bca9a2b);
sram_add_entry(0, 5, 1524, 4, 128'h4030000000000000000d94adb5f);
sram_add_entry(0, 5, 1528, 4, 128'h40300000000000000009cc28bec);
sram_add_entry(0, 5, 1532, 4, 128'h4030000000000000000f7e9401f);
sram_add_entry(0, 5, 1536, 4, 128'h4030000000000000000c81e26e4);
sram_add_entry(0, 5, 1540, 4, 128'h40300000000000000003da918ad);
sram_add_entry(0, 5, 1544, 4, 128'h403000000000000000053f821b7);
sram_add_entry(0, 5, 1548, 4, 128'h4030000000000000000e7e00d8b);
sram_add_entry(0, 5, 1552, 4, 128'h403000000000000000098e3e8fe);
sram_add_entry(0, 5, 1556, 4, 128'h4030000000000000000d66f9e32);
sram_add_entry(0, 5, 1560, 4, 128'h40300000000000000008afc2cc8);
sram_add_entry(0, 5, 1564, 4, 128'h4030000000000000000db57684a);
sram_add_entry(0, 5, 1568, 4, 128'h40300000000000000007f3dad18);
sram_add_entry(0, 5, 1572, 4, 128'h40300000000000000004a9968a9);
sram_add_entry(0, 5, 1576, 4, 128'h403000000000000000042710fa3);
sram_add_entry(0, 5, 1580, 4, 128'h40300000000000000007efb06db);
sram_add_entry(0, 5, 1584, 4, 128'h4030000000000000000958a9fd8);
sram_add_entry(0, 5, 1588, 4, 128'h40300000000000000006b82013c);
sram_add_entry(0, 5, 1592, 4, 128'h4030000000000000000eb6c6952);
sram_add_entry(0, 5, 1596, 4, 128'h4030000000000000000980df882);
sram_add_entry(0, 5, 1600, 4, 128'h403000000000000000051a3bacd);
sram_add_entry(0, 5, 1604, 4, 128'h4030000000000000000c846112e);
sram_add_entry(0, 5, 1608, 4, 128'h4030000000000000000fbb38c5d);
sram_add_entry(0, 5, 1612, 4, 128'h4030000000000000000e94cf512);
sram_add_entry(0, 5, 1616, 4, 128'h4030000000000000000ba51e5ae);
sram_add_entry(0, 5, 1620, 4, 128'h4030000000000000000202827f4);
sram_add_entry(0, 5, 1624, 4, 128'h4030000000000000000f29e4104);
sram_add_entry(0, 5, 1628, 4, 128'h40300000000000000007644bccf);
sram_add_entry(0, 5, 1632, 4, 128'h40300000000000000000dd35657);
sram_add_entry(0, 5, 1636, 4, 128'h4030000000000000000415386ed);
sram_add_entry(0, 5, 1640, 4, 128'h403000000000000000003576469);
sram_add_entry(0, 5, 1644, 4, 128'h40300000000000000001fbc279b);
sram_add_entry(0, 5, 1648, 4, 128'h4030000000000000000a271cab3);
sram_add_entry(0, 5, 1652, 4, 128'h4030000000000000000712d2a8d);
sram_add_entry(0, 5, 1656, 4, 128'h40300000000000000003fddf6b3);
sram_add_entry(0, 5, 1660, 4, 128'h40300000000000000002165be7a);
sram_add_entry(0, 5, 1664, 4, 128'h4030000000000000000448d049b);
sram_add_entry(0, 5, 1668, 4, 128'h4030000000000000000fb2d5087);
sram_add_entry(0, 5, 1672, 4, 128'h40300000000000000001e98ac81);
sram_add_entry(0, 5, 1676, 4, 128'h4030000000000000000e671ad3e);
sram_add_entry(0, 5, 1680, 4, 128'h4030000000000000000c5704dd4);
sram_add_entry(0, 5, 1684, 4, 128'h4030000000000000000b0840ac8);
sram_add_entry(0, 5, 1688, 4, 128'h4030000000000000000fa0d4b7c);
sram_add_entry(0, 5, 1692, 4, 128'h4030000000000000000ea1183e1);
sram_add_entry(0, 5, 1696, 4, 128'h4030000000000000000b91fade1);
sram_add_entry(0, 5, 1700, 4, 128'h4030000000000000000a11fde54);
sram_add_entry(0, 5, 1704, 4, 128'h403000000000000000012eff59c);
sram_add_entry(0, 5, 1708, 4, 128'h4030000000000000000db238c5d);
sram_add_entry(0, 5, 1712, 4, 128'h40300000000000000000c55954a);
sram_add_entry(0, 5, 1716, 4, 128'h40300000000000000004160f5ee);
sram_add_entry(0, 5, 1720, 4, 128'h4030000000000000000edcbd779);
sram_add_entry(0, 5, 1724, 4, 128'h4030000000000000000f4a82895);
sram_add_entry(0, 5, 1728, 4, 128'h40300000000000000001604c030);
sram_add_entry(0, 5, 1732, 4, 128'h4030000000000000000c0a439bf);
sram_add_entry(0, 5, 1736, 4, 128'h40300000000000000002a955aec);
sram_add_entry(0, 5, 1740, 4, 128'h40300000000000000002c902099);
sram_add_entry(0, 5, 1744, 4, 128'h4030000000000000000217c7717);
sram_add_entry(0, 5, 1748, 4, 128'h40300000000000000007c0ea408);
sram_add_entry(0, 5, 1752, 4, 128'h40300000000000000004d0afc5c);
sram_add_entry(0, 5, 1756, 4, 128'h4030000000000000000b8cd0eab);
sram_add_entry(0, 5, 1760, 4, 128'h4030000000000000000739e2b20);
sram_add_entry(0, 5, 1764, 4, 128'h403000000000000000034dbf565);
sram_add_entry(0, 5, 1768, 4, 128'h403000000000000000066f2d912);
sram_add_entry(0, 5, 1772, 4, 128'h4030000000000000000b7295d4e);
sram_add_entry(0, 5, 1776, 4, 128'h4030000000000000000316d5676);
sram_add_entry(0, 5, 1780, 4, 128'h403000000000000000069aa0de2);
sram_add_entry(0, 5, 1784, 4, 128'h40300000000000000007110b17d);
sram_add_entry(0, 5, 1788, 4, 128'h403000000000000000093b4e0f7);
sram_add_entry(0, 5, 1792, 4, 128'h40300000000000000004dc5b038);
sram_add_entry(0, 5, 1796, 4, 128'h4030000000000000000b9e03453);
sram_add_entry(0, 5, 1800, 4, 128'h4030000000000000000f831c057);
sram_add_entry(0, 5, 1804, 4, 128'h40300000000000000003834ff31);
sram_add_entry(0, 5, 1808, 4, 128'h4030000000000000000bcbc82bf);
sram_add_entry(0, 5, 1812, 4, 128'h40300000000000000004c1bec8b);
sram_add_entry(0, 5, 1816, 4, 128'h4030000000000000000209ec751);
sram_add_entry(0, 5, 1820, 4, 128'h40300000000000000004de18e05);
sram_add_entry(0, 5, 1824, 4, 128'h40300000000000000004f7ba449);
sram_add_entry(0, 5, 1828, 4, 128'h403000000000000000006036359);
sram_add_entry(0, 5, 1832, 4, 128'h4030000000000000000712983c2);
sram_add_entry(0, 5, 1836, 4, 128'h403000000000000000020770d60);
sram_add_entry(0, 5, 1840, 4, 128'h4030000000000000000f63206a4);
sram_add_entry(0, 5, 1844, 4, 128'h403000000000000000072a80a04);
sram_add_entry(0, 5, 1848, 4, 128'h4030000000000000000d8d85182);
sram_add_entry(0, 5, 1852, 4, 128'h4030000000000000000965e1956);
sram_add_entry(0, 5, 1856, 4, 128'h403000000000000000071bce5d1);
sram_add_entry(0, 5, 1860, 4, 128'h40300000000000000001acccf4d);
sram_add_entry(0, 5, 1864, 4, 128'h4030000000000000000be3c6600);
sram_add_entry(0, 5, 1868, 4, 128'h4030000000000000000f6b42162);
sram_add_entry(0, 5, 1872, 4, 128'h40300000000000000001ebef7e4);
sram_add_entry(0, 5, 1876, 4, 128'h4030000000000000000449b815e);
sram_add_entry(0, 5, 1880, 4, 128'h4030000000000000000f700305c);
sram_add_entry(0, 5, 1884, 4, 128'h403000000000000000071d16c63);
sram_add_entry(0, 5, 1888, 4, 128'h4030000000000000000af7769e2);
sram_add_entry(0, 5, 1892, 4, 128'h40300000000000000009238595d);
sram_add_entry(0, 5, 1896, 4, 128'h403000000000000000087abb692);
sram_add_entry(0, 5, 1900, 4, 128'h40300000000000000009f619149);
sram_add_entry(0, 5, 1904, 4, 128'h40300000000000000001c452d06);
sram_add_entry(0, 5, 1908, 4, 128'h403000000000000000047627aba);
sram_add_entry(0, 5, 1912, 4, 128'h4030000000000000000751c717c);
sram_add_entry(0, 5, 1916, 4, 128'h4030000000000000000ca65525a);
sram_add_entry(0, 5, 1920, 4, 128'h4030000000000000000b8645166);
sram_add_entry(0, 5, 1924, 4, 128'h4030000000000000000a9a978fb);
sram_add_entry(0, 5, 1928, 4, 128'h40300000000000000004f00fbb0);
sram_add_entry(0, 5, 1932, 4, 128'h4030000000000000000dc1e87e7);
sram_add_entry(0, 5, 1936, 4, 128'h40300000000000000006b81d355);
sram_add_entry(0, 5, 1940, 4, 128'h40300000000000000003e7fe58b);
sram_add_entry(0, 5, 1944, 4, 128'h4030000000000000000f3f20799);
sram_add_entry(0, 5, 1948, 4, 128'h4030000000000000000c30e1c35);
sram_add_entry(0, 5, 1952, 4, 128'h4030000000000000000da9ad8a1);
sram_add_entry(0, 5, 1956, 4, 128'h4030000000000000000fa5f7769);
sram_add_entry(0, 5, 1960, 4, 128'h4030000000000000000b1447c06);
sram_add_entry(0, 5, 1964, 4, 128'h4030000000000000000f95a7eb1);
sram_add_entry(0, 5, 1968, 4, 128'h40300000000000000009391d306);
sram_add_entry(0, 5, 1972, 4, 128'h4030000000000000000699e2b00);
sram_add_entry(0, 5, 1976, 4, 128'h4030000000000000000891868ba);
sram_add_entry(0, 5, 1980, 4, 128'h4030000000000000000a2b05c48);
sram_add_entry(0, 5, 1984, 4, 128'h4030000000000000000aac8ca5a);
sram_add_entry(0, 5, 1988, 4, 128'h40300000000000000005f8471bd);
sram_add_entry(0, 5, 1992, 4, 128'h40300000000000000000d0610bc);
sram_add_entry(0, 5, 1996, 4, 128'h403000000000000000018206fc9);
sram_add_entry(0, 5, 2000, 4, 128'h40300000000000000000ac2f36d);
sram_add_entry(0, 5, 2004, 4, 128'h403000000000000000002e748e8);
sram_add_entry(0, 5, 2008, 4, 128'h4030000000000000000f11fb9e2);
sram_add_entry(0, 5, 2012, 4, 128'h40300000000000000005b9ea50a);
sram_add_entry(0, 5, 2016, 4, 128'h4030000000000000000f227c657);
sram_add_entry(0, 5, 2020, 4, 128'h40300000000000000003515ab3b);
sram_add_entry(0, 5, 2024, 4, 128'h403000000000000000015503f8d);
sram_add_entry(0, 5, 2028, 4, 128'h403000000000000000076cc4124);
sram_add_entry(0, 5, 2032, 4, 128'h4030000000000000000d4bdec61);
sram_add_entry(0, 5, 2036, 4, 128'h4030000000000000000d2bd71db);
sram_add_entry(0, 5, 2040, 4, 128'h4030000000000000000e0a2b56f);
sram_add_entry(0, 5, 2044, 4, 128'h4030000000000000000e34d64c6);
sram_add_entry(0, 5, 2048, 4, 128'h4030000000000000000c735ad48);
sram_add_entry(0, 5, 2052, 4, 128'h40300000000000000007035214f);
sram_add_entry(0, 5, 2056, 4, 128'h4030000000000000000d2ff291a);
sram_add_entry(0, 5, 2060, 4, 128'h403000000000000000049b6cb18);
sram_add_entry(0, 5, 2064, 4, 128'h4030000000000000000c6cd4467);
sram_add_entry(0, 5, 2068, 4, 128'h4030000000000000000e90fe281);
sram_add_entry(0, 5, 2072, 4, 128'h4030000000000000000ba02a11d);
sram_add_entry(0, 5, 2076, 4, 128'h40300000000000000000253c7a3);
sram_add_entry(0, 5, 2080, 4, 128'h4030000000000000000412bb30c);
sram_add_entry(0, 5, 2084, 4, 128'h40300000000000000008d12dd56);
sram_add_entry(0, 5, 2088, 4, 128'h40300000000000000006fe0c5a1);
sram_add_entry(0, 5, 2092, 4, 128'h4030000000000000000a33b35e9);
sram_add_entry(0, 5, 2096, 4, 128'h4030000000000000000723a31b7);
sram_add_entry(0, 5, 2100, 4, 128'h40300000000000000005a350d96);
sram_add_entry(0, 5, 2104, 4, 128'h403000000000000000004006207);
sram_add_entry(0, 5, 2108, 4, 128'h4030000000000000000c702e976);
sram_add_entry(0, 5, 2112, 4, 128'h4030000000000000000b6010e92);
sram_add_entry(0, 5, 2116, 4, 128'h403000000000000000004c85212);
sram_add_entry(0, 5, 2120, 4, 128'h403000000000000000040044411);
sram_add_entry(0, 5, 2124, 4, 128'h4030000000000000000a8fb5d85);
sram_add_entry(0, 5, 2128, 4, 128'h40300000000000000004d9741f6);
sram_add_entry(0, 5, 2132, 4, 128'h4030000000000000000d3afd823);
sram_add_entry(0, 5, 2136, 4, 128'h4030000000000000000fdd6ea42);
sram_add_entry(0, 5, 2140, 4, 128'h4030000000000000000b42b3094);
sram_add_entry(0, 5, 2144, 4, 128'h40300000000000000002b35ac93);
sram_add_entry(0, 5, 2148, 4, 128'h40300000000000000001de14302);
sram_add_entry(0, 5, 2152, 4, 128'h4030000000000000000197646ab);
sram_add_entry(0, 5, 2156, 4, 128'h40300000000000000000c205d69);
sram_add_entry(0, 5, 2160, 4, 128'h40300000000000000008947a1d6);
sram_add_entry(0, 5, 2164, 4, 128'h403000000000000000006890668);
sram_add_entry(0, 5, 2168, 4, 128'h40300000000000000008bdb4cbe);
sram_add_entry(0, 5, 2172, 4, 128'h40300000000000000001969b688);
sram_add_entry(0, 5, 2176, 4, 128'h403000000000000000010e2ee9c);
sram_add_entry(0, 5, 2180, 4, 128'h4030000000000000000a7e49978);
sram_add_entry(0, 5, 2184, 4, 128'h4030000000000000000860c996f);
sram_add_entry(0, 5, 2188, 4, 128'h4030000000000000000be168c0d);
sram_add_entry(0, 5, 2192, 4, 128'h4030000000000000000f9cf89b1);
sram_add_entry(0, 5, 2196, 4, 128'h403000000000000000081261f85);
sram_add_entry(0, 5, 2200, 4, 128'h4030000000000000000e7aaa8fd);
sram_add_entry(0, 5, 2204, 4, 128'h4030000000000000000b0429c43);
sram_add_entry(0, 5, 2208, 4, 128'h40300000000000000008a4c6218);
sram_add_entry(0, 5, 2212, 4, 128'h403000000000000000095f19822);
sram_add_entry(0, 5, 2216, 4, 128'h403000000000000000045858f52);
sram_add_entry(0, 5, 2220, 4, 128'h4030000000000000000d544fa47);
sram_add_entry(0, 5, 2224, 4, 128'h4030000000000000000af1a4005);
sram_add_entry(0, 5, 2228, 4, 128'h4030000000000000000e3b732bb);
sram_add_entry(0, 5, 2232, 4, 128'h40300000000000000006194cbd6);
sram_add_entry(0, 5, 2236, 4, 128'h40300000000000000009d1b6b4b);
sram_add_entry(0, 5, 2240, 4, 128'h40300000000000000002ff0666f);
sram_add_entry(0, 5, 2244, 4, 128'h40300000000000000006913bb5f);
sram_add_entry(0, 5, 2248, 4, 128'h40300000000000000004925a9b2);
sram_add_entry(0, 5, 2252, 4, 128'h4030000000000000000cbf76125);
sram_add_entry(0, 5, 2256, 4, 128'h403000000000000000080f0a6a3);
sram_add_entry(0, 5, 2260, 4, 128'h40300000000000000001249cd1d);
sram_add_entry(0, 5, 2264, 4, 128'h4030000000000000000bc0a568e);
sram_add_entry(0, 5, 2268, 4, 128'h4030000000000000000688f87cd);
sram_add_entry(0, 5, 2272, 4, 128'h40300000000000000002960aaef);
sram_add_entry(0, 5, 2276, 4, 128'h40300000000000000005085236f);
sram_add_entry(0, 5, 2280, 4, 128'h4030000000000000000ef5d2004);
sram_add_entry(0, 5, 2284, 4, 128'h403000000000000000025b2c4aa);
sram_add_entry(0, 5, 2288, 4, 128'h4030000000000000000b972ba2f);
sram_add_entry(0, 5, 2292, 4, 128'h4030000000000000000fb315574);
sram_add_entry(0, 5, 2296, 4, 128'h40300000000000000004874d5e7);
sram_add_entry(0, 5, 2300, 4, 128'h40300000000000000008dfdecc3);
sram_add_entry(0, 5, 2304, 4, 128'h4030000000000000000cce699ec);
sram_add_entry(0, 5, 2308, 4, 128'h4030000000000000000785b1a49);
sram_add_entry(0, 5, 2312, 4, 128'h4030000000000000000ebe00791);
sram_add_entry(0, 5, 2316, 4, 128'h4030000000000000000c3beb879);
sram_add_entry(0, 5, 2320, 4, 128'h4030000000000000000e4c31860);
sram_add_entry(0, 5, 2324, 4, 128'h40300000000000000000d6fbba7);
sram_add_entry(0, 5, 2328, 4, 128'h4030000000000000000f165457d);
sram_add_entry(0, 5, 2332, 4, 128'h40300000000000000003805f41d);
sram_add_entry(0, 5, 2336, 4, 128'h403000000000000000058045c79);
sram_add_entry(0, 5, 2340, 4, 128'h4030000000000000000b77beed9);
sram_add_entry(0, 5, 2344, 4, 128'h4030000000000000000364e16c5);
sram_add_entry(0, 5, 2348, 4, 128'h4030000000000000000379023ab);
sram_add_entry(0, 5, 2352, 4, 128'h40300000000000000001f3f2a95);
sram_add_entry(0, 5, 2356, 4, 128'h40300000000000000006317bf23);
sram_add_entry(0, 5, 2360, 4, 128'h403000000000000000075d392b5);
sram_add_entry(0, 5, 2364, 4, 128'h4030000000000000000d7f4bb13);
sram_add_entry(0, 5, 2368, 4, 128'h4030000000000000000bdf1b95a);
sram_add_entry(0, 5, 2372, 4, 128'h4030000000000000000ff3fdc47);
sram_add_entry(0, 5, 2376, 4, 128'h4030000000000000000fe817339);
sram_add_entry(0, 5, 2380, 4, 128'h4030000000000000000b670bd6a);
sram_add_entry(0, 5, 2384, 4, 128'h403000000000000000080fb1afb);
sram_add_entry(0, 5, 2388, 4, 128'h40300000000000000007e488471);
sram_add_entry(0, 5, 2392, 4, 128'h4030000000000000000180ab825);
sram_add_entry(0, 5, 2396, 4, 128'h4030000000000000000432afc9f);
sram_add_entry(0, 5, 2400, 4, 128'h40300000000000000000e23107c);
sram_add_entry(0, 5, 2404, 4, 128'h4030000000000000000266062f1);
sram_add_entry(0, 5, 2408, 4, 128'h40300000000000000002ff8a855);
sram_add_entry(0, 5, 2412, 4, 128'h40300000000000000001ba59a2e);
sram_add_entry(0, 5, 2416, 4, 128'h40300000000000000003a0d39c7);
sram_add_entry(0, 5, 2420, 4, 128'h403000000000000000098c7b823);
sram_add_entry(0, 5, 2424, 4, 128'h40300000000000000005462a053);
sram_add_entry(0, 5, 2428, 4, 128'h4030000000000000000ced324b2);
sram_add_entry(0, 5, 2432, 4, 128'h40300000000000000007808026c);
sram_add_entry(0, 5, 2436, 4, 128'h403000000000000000076544554);
sram_add_entry(0, 5, 2440, 4, 128'h4030000000000000000587748f1);
sram_add_entry(0, 5, 2444, 4, 128'h4030000000000000000f759b497);
sram_add_entry(0, 5, 2448, 4, 128'h403000000000000000049dd7a37);
sram_add_entry(0, 5, 2452, 4, 128'h4030000000000000000b16968b0);
sram_add_entry(0, 5, 2456, 4, 128'h403000000000000000080c27aff);
sram_add_entry(0, 5, 2460, 4, 128'h4030000000000000000d5249c05);
sram_add_entry(0, 5, 2464, 4, 128'h40300000000000000009b3bb04a);
sram_add_entry(0, 5, 2468, 4, 128'h4030000000000000000c4f06715);
sram_add_entry(0, 5, 2472, 4, 128'h403000000000000000060e58984);
sram_add_entry(0, 5, 2476, 4, 128'h4030000000000000000a69c4dec);
sram_add_entry(0, 5, 2480, 4, 128'h40300000000000000009996b95e);
sram_add_entry(0, 5, 2484, 4, 128'h4030000000000000000b3533b00);
sram_add_entry(0, 5, 2488, 4, 128'h40300000000000000006034dd18);
sram_add_entry(0, 5, 2492, 4, 128'h403000000000000000074e86cc8);
sram_add_entry(0, 5, 2496, 4, 128'h4030000000000000000a06c8f64);
sram_add_entry(0, 5, 2500, 4, 128'h40300000000000000003f2bc9a0);
sram_add_entry(0, 5, 2504, 4, 128'h4030000000000000000f81585e9);
sram_add_entry(0, 5, 2508, 4, 128'h403000000000000000097515402);
sram_add_entry(0, 5, 2512, 4, 128'h403000000000000000002a07f05);
sram_add_entry(0, 5, 2516, 4, 128'h40300000000000000002bc32216);
sram_add_entry(0, 5, 2520, 4, 128'h4030000000000000000909c5b0d);
sram_add_entry(0, 5, 2524, 4, 128'h4030000000000000000e5dcf0e6);
sram_add_entry(0, 5, 2528, 4, 128'h4030000000000000000965ce467);
sram_add_entry(0, 5, 2532, 4, 128'h40300000000000000002fe7f356);
sram_add_entry(0, 5, 2536, 4, 128'h403000000000000000030d25e12);
sram_add_entry(0, 5, 2540, 4, 128'h40300000000000000004bb8ac18);
sram_add_entry(0, 5, 2544, 4, 128'h403000000000000000044f4a58a);
sram_add_entry(0, 5, 2548, 4, 128'h40300000000000000000f501287);
sram_add_entry(0, 5, 2552, 4, 128'h40300000000000000007eaf6d4f);
sram_add_entry(0, 5, 2556, 4, 128'h4030000000000000000d82212f1);
sram_add_entry(0, 5, 2560, 4, 128'h4030000000000000000ec1625ea);
sram_add_entry(0, 5, 2564, 4, 128'h403000000000000000074cae5e1);
sram_add_entry(0, 5, 2568, 4, 128'h40300000000000000001fe03adc);
sram_add_entry(0, 5, 2572, 4, 128'h4030000000000000000e0ce0e82);
sram_add_entry(0, 5, 2576, 4, 128'h40300000000000000005f82b623);
sram_add_entry(0, 5, 2580, 4, 128'h403000000000000000007e2be26);
sram_add_entry(0, 5, 2584, 4, 128'h4030000000000000000b4c4d344);
sram_add_entry(0, 5, 2588, 4, 128'h403000000000000000002ecd929);
sram_add_entry(0, 5, 2592, 4, 128'h4030000000000000000c583cf7b);
sram_add_entry(0, 5, 2596, 4, 128'h4030000000000000000f4373181);
sram_add_entry(0, 5, 2600, 4, 128'h4030000000000000000c69ba9fb);
sram_add_entry(0, 5, 2604, 4, 128'h40300000000000000008b43e12f);
sram_add_entry(0, 5, 2608, 4, 128'h40300000000000000001a7a8797);
sram_add_entry(0, 5, 2612, 4, 128'h40300000000000000006dcbaa62);
sram_add_entry(0, 5, 2616, 4, 128'h4030000000000000000046285e0);
sram_add_entry(0, 5, 2620, 4, 128'h4030000000000000000c9e05443);
sram_add_entry(0, 5, 2624, 4, 128'h40300000000000000007f136176);
sram_add_entry(0, 5, 2628, 4, 128'h40300000000000000000a9a396f);
sram_add_entry(0, 5, 2632, 4, 128'h4030000000000000000d535e00d);
sram_add_entry(0, 5, 2636, 4, 128'h403000000000000000076394b0c);
sram_add_entry(0, 5, 2640, 4, 128'h40300000000000000000a330561);
sram_add_entry(0, 5, 2644, 4, 128'h403000000000000000043b01a49);
sram_add_entry(0, 5, 2648, 4, 128'h4030000000000000000ff999355);
sram_add_entry(0, 5, 2652, 4, 128'h4030000000000000000a5eddcfb);
sram_add_entry(0, 5, 2656, 4, 128'h403000000000000000045f82b33);
sram_add_entry(0, 5, 2660, 4, 128'h40300000000000000004a4c1e12);
sram_add_entry(0, 5, 2664, 4, 128'h40300000000000000003b8a6857);
sram_add_entry(0, 5, 2668, 4, 128'h4030000000000000000b1e16a4c);
sram_add_entry(0, 5, 2672, 4, 128'h4030000000000000000fce324ac);
sram_add_entry(0, 5, 2676, 4, 128'h4030000000000000000e619bc20);
sram_add_entry(0, 5, 2680, 4, 128'h40300000000000000002caded6b);
sram_add_entry(0, 5, 2684, 4, 128'h40300000000000000003b50576b);
sram_add_entry(0, 5, 2688, 4, 128'h4030000000000000000640ef1ce);
sram_add_entry(0, 5, 2692, 4, 128'h4030000000000000000f21564b1);
sram_add_entry(0, 5, 2696, 4, 128'h403000000000000000025f779da);
sram_add_entry(0, 5, 2700, 4, 128'h4030000000000000000425844e1);
sram_add_entry(0, 5, 2704, 4, 128'h4030000000000000000e8c91e81);
sram_add_entry(0, 5, 2708, 4, 128'h40300000000000000008c9c6fa7);
sram_add_entry(0, 5, 2712, 4, 128'h403000000000000000079a69237);
sram_add_entry(0, 5, 2716, 4, 128'h40300000000000000001db22a87);
sram_add_entry(0, 5, 2720, 4, 128'h4030000000000000000243c5486);
sram_add_entry(0, 5, 2724, 4, 128'h4030000000000000000935fc3ce);
sram_add_entry(0, 5, 2728, 4, 128'h4030000000000000000590e4270);
sram_add_entry(0, 5, 2732, 4, 128'h4030000000000000000707e28f6);
sram_add_entry(0, 5, 2736, 4, 128'h4030000000000000000dae57a3d);
sram_add_entry(0, 5, 2740, 4, 128'h4030000000000000000b87638d9);
sram_add_entry(0, 5, 2744, 4, 128'h4030000000000000000d4807ce9);
sram_add_entry(0, 5, 2748, 4, 128'h40300000000000000008c9c8a90);
sram_add_entry(0, 5, 2752, 4, 128'h4030000000000000000785a9702);
sram_add_entry(0, 5, 2756, 4, 128'h4030000000000000000b1259e5a);
sram_add_entry(0, 5, 2760, 4, 128'h40300000000000000009cb6c8e9);
sram_add_entry(0, 5, 2764, 4, 128'h4030000000000000000641e0603);
sram_add_entry(0, 5, 2768, 4, 128'h4030000000000000000fa391441);
sram_add_entry(0, 5, 2772, 4, 128'h40300000000000000002b6458e0);
sram_add_entry(0, 5, 2776, 4, 128'h4030000000000000000268cf6b2);
sram_add_entry(0, 5, 2780, 4, 128'h40300000000000000007858cb29);
sram_add_entry(0, 5, 2784, 4, 128'h4030000000000000000c0447d97);
sram_add_entry(0, 5, 2788, 4, 128'h40300000000000000000abd5331);
sram_add_entry(0, 5, 2792, 4, 128'h40300000000000000008ccb7b91);
sram_add_entry(0, 5, 2796, 4, 128'h4030000000000000000722790a4);
sram_add_entry(0, 5, 2800, 4, 128'h403000000000000000001de04b8);
sram_add_entry(0, 6, 0, 4, 128'h7ab000000000000000000deadbf);
sram_add_entry(0, 6, 4, 4, 128'h40300000000000000000000ec67);
sram_add_entry(0, 6, 8, 4, 128'h40300000000000000000000ca33);
sram_add_entry(0, 6, 12, 4, 128'h403000000000000000000006d67);
sram_add_entry(0, 6, 16, 4, 128'h40300000000000000000000c411);
sram_add_entry(0, 6, 20, 4, 128'h40300000000000000000000e871);
sram_add_entry(0, 6, 24, 4, 128'h40300000000000000000000434d);
sram_add_entry(0, 6, 28, 4, 128'h40300000000000000000000bc90);
sram_add_entry(0, 6, 32, 4, 128'h403000000000000000000003182);
sram_add_entry(0, 6, 36, 4, 128'h40300000000000000000000f995);
sram_add_entry(0, 6, 40, 4, 128'h40300000000000000000000ab9b);
sram_add_entry(0, 6, 44, 4, 128'h403000000000000000000003f0e);
sram_add_entry(0, 6, 48, 4, 128'h403000000000000000000000a49);
sram_add_entry(0, 6, 52, 4, 128'h403000000000000000000009ced);
sram_add_entry(0, 6, 56, 4, 128'h40300000000000000000000fa16);
sram_add_entry(0, 6, 60, 4, 128'h403000000000000000000000bf3);
sram_add_entry(0, 6, 64, 4, 128'h40300000000000000000000ecf9);
sram_add_entry(0, 6, 68, 4, 128'h40300000000000000000000273b);
sram_add_entry(0, 6, 72, 4, 128'h403000000000000000000007d62);
sram_add_entry(0, 6, 76, 4, 128'h403000000000000000000003658);
sram_add_entry(0, 6, 80, 4, 128'h40300000000000000000000d34c);
sram_add_entry(0, 6, 84, 4, 128'h40300000000000000000000a11e);
sram_add_entry(0, 6, 88, 4, 128'h40300000000000000000000cdb1);
sram_add_entry(0, 6, 92, 4, 128'h40300000000000000000000cb23);
sram_add_entry(0, 6, 96, 4, 128'h403000000000000000000004f15);
sram_add_entry(0, 6, 100, 4, 128'h4030000000000000000000000f6);
sram_add_entry(0, 6, 104, 4, 128'h403000000000000000000008a2b);
sram_add_entry(0, 6, 108, 4, 128'h403000000000000000000000b21);
sram_add_entry(0, 6, 112, 4, 128'h403000000000000000000001699);
sram_add_entry(0, 6, 116, 4, 128'h4030000000000000000000001d0);
sram_add_entry(0, 6, 120, 4, 128'h40300000000000000000000daf2);
sram_add_entry(0, 6, 124, 4, 128'h40300000000000000000000317c);
sram_add_entry(0, 6, 128, 4, 128'h403000000000000000000005312);
sram_add_entry(0, 6, 132, 4, 128'h40300000000000000000000cd1a);
sram_add_entry(0, 6, 136, 4, 128'h4030000000000000000000024e6);
sram_add_entry(0, 6, 140, 4, 128'h403000000000000000000008650);
sram_add_entry(0, 6, 144, 4, 128'h40300000000000000000000948a);
sram_add_entry(0, 6, 148, 4, 128'h403000000000000000000003b16);
sram_add_entry(0, 6, 152, 4, 128'h40300000000000000000000d1cc);
sram_add_entry(0, 6, 156, 4, 128'h40300000000000000000000ed39);
sram_add_entry(0, 6, 160, 4, 128'h403000000000000000000004552);
sram_add_entry(0, 6, 164, 4, 128'h403000000000000000000003604);
sram_add_entry(0, 6, 168, 4, 128'h40300000000000000000000128b);
sram_add_entry(0, 6, 172, 4, 128'h40300000000000000000000e052);
sram_add_entry(0, 6, 176, 4, 128'h403000000000000000000009626);
sram_add_entry(0, 6, 180, 4, 128'h403000000000000000000006ae6);
sram_add_entry(0, 6, 184, 4, 128'h403000000000000000000005c87);
sram_add_entry(0, 6, 188, 4, 128'h403000000000000000000008b78);
sram_add_entry(0, 6, 192, 4, 128'h403000000000000000000004875);
sram_add_entry(0, 6, 196, 4, 128'h403000000000000000000002d1e);
sram_add_entry(0, 6, 200, 4, 128'h403000000000000000000005b49);
sram_add_entry(0, 6, 204, 4, 128'h4030000000000000000000059b7);
sram_add_entry(0, 6, 208, 4, 128'h40300000000000000000000e851);
sram_add_entry(0, 6, 212, 4, 128'h403000000000000000000005ca1);
sram_add_entry(0, 6, 216, 4, 128'h403000000000000000000007ba3);
sram_add_entry(0, 6, 220, 4, 128'h4030000000000000000000002c4);
sram_add_entry(0, 6, 224, 4, 128'h403000000000000000000004df4);
sram_add_entry(0, 6, 228, 4, 128'h403000000000000000000006933);
sram_add_entry(0, 6, 232, 4, 128'h40300000000000000000000e4f4);
sram_add_entry(0, 6, 236, 4, 128'h40300000000000000000000e474);
sram_add_entry(0, 6, 240, 4, 128'h40300000000000000000000b8d7);
sram_add_entry(0, 6, 244, 4, 128'h403000000000000000000003227);
sram_add_entry(0, 6, 248, 4, 128'h40300000000000000000000aae6);
sram_add_entry(0, 6, 252, 4, 128'h4030000000000000000000062c4);
sram_add_entry(0, 6, 256, 4, 128'h40300000000000000000000dd68);
sram_add_entry(0, 6, 260, 4, 128'h403000000000000000000007e73);
sram_add_entry(0, 6, 264, 4, 128'h4030000000000000000000003af);
sram_add_entry(0, 6, 268, 4, 128'h4030000000000000000000048de);
sram_add_entry(0, 6, 272, 4, 128'h403000000000000000000000efd);
sram_add_entry(0, 6, 276, 4, 128'h40300000000000000000000e419);
sram_add_entry(0, 6, 280, 4, 128'h403000000000000000000009356);
sram_add_entry(0, 6, 284, 4, 128'h40300000000000000000000a8b9);
sram_add_entry(0, 6, 288, 4, 128'h4030000000000000000000064c1);
sram_add_entry(0, 6, 292, 4, 128'h40300000000000000000000b6da);
sram_add_entry(0, 6, 296, 4, 128'h40300000000000000000000ea32);
sram_add_entry(0, 6, 300, 4, 128'h403000000000000000000005eed);
sram_add_entry(0, 6, 304, 4, 128'h40300000000000000000000faf4);
sram_add_entry(0, 6, 308, 4, 128'h403000000000000000000007a2c);
sram_add_entry(0, 6, 312, 4, 128'h40300000000000000000000f957);
sram_add_entry(0, 6, 316, 4, 128'h403000000000000000000005b6b);
sram_add_entry(0, 6, 320, 4, 128'h403000000000000000000003d98);
sram_add_entry(0, 6, 324, 4, 128'h40300000000000000000000f6bf);
sram_add_entry(0, 6, 328, 4, 128'h40300000000000000000000933e);
sram_add_entry(0, 6, 332, 4, 128'h403000000000000000000004e1f);
sram_add_entry(0, 6, 336, 4, 128'h403000000000000000000007a3d);
sram_add_entry(0, 6, 340, 4, 128'h403000000000000000000007d64);
sram_add_entry(0, 6, 344, 4, 128'h40300000000000000000000dfa6);
sram_add_entry(0, 6, 348, 4, 128'h40300000000000000000000e19a);
sram_add_entry(0, 6, 352, 4, 128'h4030000000000000000000066d1);
sram_add_entry(0, 6, 356, 4, 128'h40300000000000000000000f6c4);
sram_add_entry(0, 6, 360, 4, 128'h40300000000000000000000acc9);
sram_add_entry(0, 6, 364, 4, 128'h40300000000000000000000a5aa);
sram_add_entry(0, 6, 368, 4, 128'h40300000000000000000000777f);
sram_add_entry(0, 6, 372, 4, 128'h40300000000000000000000f0f0);
sram_add_entry(0, 6, 376, 4, 128'h40300000000000000000000cfbb);
sram_add_entry(0, 6, 380, 4, 128'h403000000000000000000002c19);
sram_add_entry(0, 6, 384, 4, 128'h4030000000000000000000024d4);
sram_add_entry(0, 6, 388, 4, 128'h403000000000000000000005ffc);
sram_add_entry(0, 6, 392, 4, 128'h40300000000000000000000acf5);
sram_add_entry(0, 6, 396, 4, 128'h40300000000000000000000894c);
sram_add_entry(0, 6, 400, 4, 128'h4030000000000000000000017ab);
sram_add_entry(0, 6, 404, 4, 128'h403000000000000000000001075);
sram_add_entry(0, 6, 408, 4, 128'h403000000000000000000005677);
sram_add_entry(0, 6, 412, 4, 128'h403000000000000000000001b39);
sram_add_entry(0, 6, 416, 4, 128'h403000000000000000000003a80);
sram_add_entry(0, 6, 420, 4, 128'h403000000000000000000003017);
sram_add_entry(0, 6, 424, 4, 128'h403000000000000000000009202);
sram_add_entry(0, 6, 428, 4, 128'h4030000000000000000000074cd);
sram_add_entry(0, 6, 432, 4, 128'h403000000000000000000005c5f);
sram_add_entry(0, 6, 436, 4, 128'h403000000000000000000001117);
sram_add_entry(0, 6, 440, 4, 128'h40300000000000000000000e794);
sram_add_entry(0, 6, 444, 4, 128'h40300000000000000000000a456);
sram_add_entry(0, 6, 448, 4, 128'h40300000000000000000000cfdd);
sram_add_entry(0, 6, 452, 4, 128'h40300000000000000000000d835);
sram_add_entry(0, 6, 456, 4, 128'h40300000000000000000000dd49);
sram_add_entry(0, 6, 460, 4, 128'h403000000000000000000007570);
sram_add_entry(0, 6, 464, 4, 128'h40300000000000000000000b255);
sram_add_entry(0, 6, 468, 4, 128'h403000000000000000000006980);
sram_add_entry(0, 6, 472, 4, 128'h403000000000000000000008260);
sram_add_entry(0, 6, 476, 4, 128'h40300000000000000000000a205);
sram_add_entry(0, 6, 480, 4, 128'h40300000000000000000000304d);
sram_add_entry(0, 6, 484, 4, 128'h40300000000000000000000fb08);
sram_add_entry(0, 6, 488, 4, 128'h40300000000000000000000fa71);
sram_add_entry(0, 6, 492, 4, 128'h40300000000000000000000e4d8);
sram_add_entry(0, 6, 496, 4, 128'h403000000000000000000001c3e);
sram_add_entry(0, 6, 500, 4, 128'h403000000000000000000004931);
sram_add_entry(0, 6, 504, 4, 128'h4030000000000000000000084b5);
sram_add_entry(0, 6, 508, 4, 128'h403000000000000000000000711);
sram_add_entry(0, 6, 512, 4, 128'h40300000000000000000000ca64);
sram_add_entry(0, 6, 516, 4, 128'h40300000000000000000000d669);
sram_add_entry(0, 6, 520, 4, 128'h403000000000000000000004363);
sram_add_entry(0, 6, 524, 4, 128'h40300000000000000000000f838);
sram_add_entry(0, 6, 528, 4, 128'h403000000000000000000008a28);
sram_add_entry(0, 6, 532, 4, 128'h40300000000000000000000811a);
sram_add_entry(0, 6, 536, 4, 128'h40300000000000000000000040c);
sram_add_entry(0, 6, 540, 4, 128'h4030000000000000000000041ac);
sram_add_entry(0, 6, 544, 4, 128'h403000000000000000000004b1b);
sram_add_entry(0, 6, 548, 4, 128'h40300000000000000000000b214);
sram_add_entry(0, 6, 552, 4, 128'h40300000000000000000000504f);
sram_add_entry(0, 6, 556, 4, 128'h40300000000000000000000ae5d);
sram_add_entry(0, 6, 560, 4, 128'h40300000000000000000000914b);
sram_add_entry(0, 6, 564, 4, 128'h403000000000000000000004c67);
sram_add_entry(0, 6, 568, 4, 128'h4030000000000000000000025f9);
sram_add_entry(0, 6, 572, 4, 128'h403000000000000000000002323);
sram_add_entry(0, 6, 576, 4, 128'h403000000000000000000003f89);
sram_add_entry(0, 6, 580, 4, 128'h4030000000000000000000005c3);
sram_add_entry(0, 6, 584, 4, 128'h403000000000000000000008362);
sram_add_entry(0, 6, 588, 4, 128'h40300000000000000000000d4ed);
sram_add_entry(0, 6, 592, 4, 128'h403000000000000000000001634);
sram_add_entry(0, 6, 596, 4, 128'h403000000000000000000006bb4);
sram_add_entry(0, 6, 600, 4, 128'h403000000000000000000008ca3);
sram_add_entry(0, 6, 604, 4, 128'h40300000000000000000000c978);
sram_add_entry(0, 6, 608, 4, 128'h40300000000000000000000f216);
sram_add_entry(0, 6, 612, 4, 128'h40300000000000000000000cd29);
sram_add_entry(0, 6, 616, 4, 128'h403000000000000000000005114);
sram_add_entry(0, 6, 620, 4, 128'h403000000000000000000005ffc);
sram_add_entry(0, 6, 624, 4, 128'h40300000000000000000000efa8);
sram_add_entry(0, 6, 628, 4, 128'h4030000000000000000000000a3);
sram_add_entry(0, 6, 632, 4, 128'h403000000000000000000005bcb);
sram_add_entry(0, 6, 636, 4, 128'h4030000000000000000000034d2);
sram_add_entry(0, 6, 640, 4, 128'h40300000000000000000000b6ed);
sram_add_entry(0, 6, 644, 4, 128'h403000000000000000000002d7a);
sram_add_entry(0, 6, 648, 4, 128'h4030000000000000000000053b8);
sram_add_entry(0, 6, 652, 4, 128'h403000000000000000000009151);
sram_add_entry(0, 6, 656, 4, 128'h403000000000000000000008bc6);
sram_add_entry(0, 6, 660, 4, 128'h4030000000000000000000074ce);
sram_add_entry(0, 6, 664, 4, 128'h40300000000000000000000300e);
sram_add_entry(0, 6, 668, 4, 128'h403000000000000000000006347);
sram_add_entry(0, 6, 672, 4, 128'h403000000000000000000008a2f);
sram_add_entry(0, 6, 676, 4, 128'h40300000000000000000000775b);
sram_add_entry(0, 6, 680, 4, 128'h40300000000000000000000b202);
sram_add_entry(0, 6, 684, 4, 128'h4030000000000000000000043c7);
sram_add_entry(0, 6, 688, 4, 128'h4030000000000000000000077bb);
sram_add_entry(0, 6, 692, 4, 128'h40300000000000000000000567e);
sram_add_entry(0, 6, 696, 4, 128'h403000000000000000000008d37);
sram_add_entry(0, 6, 700, 4, 128'h40300000000000000000000f369);
sram_add_entry(0, 6, 704, 4, 128'h403000000000000000000003a0f);
sram_add_entry(0, 6, 708, 4, 128'h40300000000000000000000a1f5);
sram_add_entry(0, 6, 712, 4, 128'h4030000000000000000000076a9);
sram_add_entry(0, 6, 716, 4, 128'h403000000000000000000001474);
sram_add_entry(0, 6, 720, 4, 128'h4030000000000000000000052e6);
sram_add_entry(0, 6, 724, 4, 128'h403000000000000000000002f51);
sram_add_entry(0, 6, 728, 4, 128'h40300000000000000000000652b);
sram_add_entry(0, 6, 732, 4, 128'h40300000000000000000000e3f9);
sram_add_entry(0, 6, 736, 4, 128'h403000000000000000000000a7a);
sram_add_entry(0, 6, 740, 4, 128'h40300000000000000000000b249);
sram_add_entry(0, 6, 744, 4, 128'h4030000000000000000000032a0);
sram_add_entry(0, 6, 748, 4, 128'h403000000000000000000006074);
sram_add_entry(0, 6, 752, 4, 128'h403000000000000000000003737);
sram_add_entry(0, 6, 756, 4, 128'h403000000000000000000002dfa);
sram_add_entry(0, 6, 760, 4, 128'h40300000000000000000000a1f2);
sram_add_entry(0, 6, 764, 4, 128'h403000000000000000000004653);
sram_add_entry(0, 6, 768, 4, 128'h4030000000000000000000027fb);
sram_add_entry(0, 6, 772, 4, 128'h40300000000000000000000e2cf);
sram_add_entry(0, 6, 776, 4, 128'h40300000000000000000000c65c);
sram_add_entry(0, 6, 780, 4, 128'h40300000000000000000000cfb9);
sram_add_entry(0, 6, 784, 4, 128'h403000000000000000000000295);
sram_add_entry(0, 6, 788, 4, 128'h40300000000000000000000639d);
sram_add_entry(0, 6, 792, 4, 128'h403000000000000000000007807);
sram_add_entry(0, 6, 796, 4, 128'h4030000000000000000000014ab);
sram_add_entry(0, 6, 800, 4, 128'h403000000000000000000002540);
sram_add_entry(0, 6, 804, 4, 128'h40300000000000000000000a6b5);
sram_add_entry(0, 6, 808, 4, 128'h40300000000000000000000349d);
sram_add_entry(0, 6, 812, 4, 128'h40300000000000000000000d281);
sram_add_entry(0, 6, 816, 4, 128'h40300000000000000000000142d);
sram_add_entry(0, 6, 820, 4, 128'h403000000000000000000006d0d);
sram_add_entry(0, 6, 824, 4, 128'h40300000000000000000000e636);
sram_add_entry(0, 6, 828, 4, 128'h40300000000000000000000a342);
sram_add_entry(0, 6, 832, 4, 128'h4030000000000000000000025d3);
sram_add_entry(0, 6, 836, 4, 128'h403000000000000000000000acf);
sram_add_entry(0, 6, 840, 4, 128'h4030000000000000000000058ca);
sram_add_entry(0, 6, 844, 4, 128'h40300000000000000000000b00e);
sram_add_entry(0, 6, 848, 4, 128'h40300000000000000000000b9c1);
sram_add_entry(0, 6, 852, 4, 128'h40300000000000000000000091d);
sram_add_entry(0, 6, 856, 4, 128'h403000000000000000000008e15);
sram_add_entry(0, 6, 860, 4, 128'h40300000000000000000000ff14);
sram_add_entry(0, 6, 864, 4, 128'h4030000000000000000000057fa);
sram_add_entry(0, 6, 868, 4, 128'h40300000000000000000000da3f);
sram_add_entry(0, 6, 872, 4, 128'h403000000000000000000000f47);
sram_add_entry(0, 6, 876, 4, 128'h40300000000000000000000ad05);
sram_add_entry(0, 6, 880, 4, 128'h403000000000000000000005563);
sram_add_entry(0, 6, 884, 4, 128'h40300000000000000000000534f);
sram_add_entry(0, 6, 888, 4, 128'h40300000000000000000000327f);
sram_add_entry(0, 6, 892, 4, 128'h403000000000000000000007e5b);
sram_add_entry(0, 6, 896, 4, 128'h40300000000000000000000adda);
sram_add_entry(0, 6, 900, 4, 128'h40300000000000000000000c981);
sram_add_entry(0, 6, 904, 4, 128'h40300000000000000000000d139);
sram_add_entry(0, 6, 908, 4, 128'h403000000000000000000002513);
sram_add_entry(0, 6, 912, 4, 128'h40300000000000000000000327d);
sram_add_entry(0, 6, 916, 4, 128'h403000000000000000000009e05);
sram_add_entry(0, 6, 920, 4, 128'h40300000000000000000000f241);
sram_add_entry(0, 6, 924, 4, 128'h403000000000000000000001dee);
sram_add_entry(0, 6, 928, 4, 128'h40300000000000000000000d55e);
sram_add_entry(0, 6, 932, 4, 128'h4030000000000000000000025de);
sram_add_entry(0, 6, 936, 4, 128'h40300000000000000000000df66);
sram_add_entry(0, 6, 940, 4, 128'h40300000000000000000000260e);
sram_add_entry(0, 6, 944, 4, 128'h4030000000000000000000011f9);
sram_add_entry(0, 6, 948, 4, 128'h403000000000000000000007851);
sram_add_entry(0, 6, 952, 4, 128'h403000000000000000000004bb5);
sram_add_entry(0, 6, 956, 4, 128'h4030000000000000000000058ad);
sram_add_entry(0, 6, 960, 4, 128'h40300000000000000000000cd39);
sram_add_entry(0, 6, 964, 4, 128'h403000000000000000000004594);
sram_add_entry(0, 6, 968, 4, 128'h403000000000000000000009e8b);
sram_add_entry(0, 6, 972, 4, 128'h403000000000000000000007e25);
sram_add_entry(0, 6, 976, 4, 128'h403000000000000000000009c66);
sram_add_entry(0, 6, 980, 4, 128'h40300000000000000000000067e);
sram_add_entry(0, 6, 984, 4, 128'h403000000000000000000001f05);
sram_add_entry(0, 6, 988, 4, 128'h403000000000000000000003663);
sram_add_entry(0, 6, 992, 4, 128'h40300000000000000000000c3fb);
sram_add_entry(0, 6, 996, 4, 128'h40300000000000000000000689d);
sram_add_entry(0, 6, 1000, 4, 128'h403000000000000000000006519);
sram_add_entry(0, 6, 1004, 4, 128'h40300000000000000000000efd8);
sram_add_entry(0, 6, 1008, 4, 128'h40300000000000000000000cf65);
sram_add_entry(0, 6, 1012, 4, 128'h403000000000000000000002090);
sram_add_entry(0, 6, 1016, 4, 128'h403000000000000000000007423);
sram_add_entry(0, 6, 1020, 4, 128'h403000000000000000000002ac0);
sram_add_entry(0, 6, 1024, 4, 128'h403000000000000000000005ce1);
sram_add_entry(0, 6, 1028, 4, 128'h403000000000000000000002f49);
sram_add_entry(0, 6, 1032, 4, 128'h40300000000000000000000e74d);
sram_add_entry(0, 6, 1036, 4, 128'h40300000000000000000000fe3a);
sram_add_entry(0, 6, 1040, 4, 128'h403000000000000000000001570);
sram_add_entry(0, 6, 1044, 4, 128'h4030000000000000000000096ed);
sram_add_entry(0, 6, 1048, 4, 128'h403000000000000000000002b86);
sram_add_entry(0, 6, 1052, 4, 128'h4030000000000000000000003c2);
sram_add_entry(0, 6, 1056, 4, 128'h40300000000000000000000d542);
sram_add_entry(0, 6, 1060, 4, 128'h403000000000000000000005df5);
sram_add_entry(0, 6, 1064, 4, 128'h403000000000000000000008aa0);
sram_add_entry(0, 6, 1068, 4, 128'h40300000000000000000000a9a3);
sram_add_entry(0, 6, 1072, 4, 128'h4030000000000000000000042d3);
sram_add_entry(0, 6, 1076, 4, 128'h403000000000000000000008837);
sram_add_entry(0, 6, 1080, 4, 128'h403000000000000000000003ced);
sram_add_entry(0, 6, 1084, 4, 128'h4030000000000000000000048b0);
sram_add_entry(0, 6, 1088, 4, 128'h403000000000000000000000d5f);
sram_add_entry(0, 6, 1092, 4, 128'h40300000000000000000000f9fd);
sram_add_entry(0, 6, 1096, 4, 128'h4030000000000000000000012ac);
sram_add_entry(0, 6, 1100, 4, 128'h403000000000000000000009222);
sram_add_entry(0, 6, 1104, 4, 128'h403000000000000000000004182);
sram_add_entry(0, 6, 1108, 4, 128'h403000000000000000000009201);
sram_add_entry(0, 6, 1112, 4, 128'h403000000000000000000009c52);
sram_add_entry(0, 6, 1116, 4, 128'h403000000000000000000008583);
sram_add_entry(0, 6, 1120, 4, 128'h40300000000000000000000f1e2);
sram_add_entry(0, 6, 1124, 4, 128'h40300000000000000000000b68d);
sram_add_entry(0, 6, 1128, 4, 128'h4030000000000000000000022c5);
sram_add_entry(0, 6, 1132, 4, 128'h4030000000000000000000035a0);
sram_add_entry(0, 6, 1136, 4, 128'h40300000000000000000000d202);
sram_add_entry(0, 6, 1140, 4, 128'h4030000000000000000000087af);
sram_add_entry(0, 6, 1144, 4, 128'h40300000000000000000000f3b0);
sram_add_entry(0, 6, 1148, 4, 128'h40300000000000000000000646e);
sram_add_entry(0, 6, 1152, 4, 128'h40300000000000000000000227e);
sram_add_entry(0, 6, 1156, 4, 128'h40300000000000000000000dbb4);
sram_add_entry(0, 6, 1160, 4, 128'h403000000000000000000002830);
sram_add_entry(0, 6, 1164, 4, 128'h403000000000000000000000f47);
sram_add_entry(0, 6, 1168, 4, 128'h403000000000000000000006e3a);
sram_add_entry(0, 6, 1172, 4, 128'h4030000000000000000000013f3);
sram_add_entry(0, 6, 1176, 4, 128'h403000000000000000000004667);
sram_add_entry(0, 6, 1180, 4, 128'h4030000000000000000000039b8);
sram_add_entry(0, 6, 1184, 4, 128'h4030000000000000000000054e5);
sram_add_entry(0, 6, 1188, 4, 128'h4030000000000000000000058ec);
sram_add_entry(0, 6, 1192, 4, 128'h403000000000000000000006869);
sram_add_entry(0, 6, 1196, 4, 128'h403000000000000000000006bbe);
sram_add_entry(0, 6, 1200, 4, 128'h403000000000000000000007815);
sram_add_entry(0, 6, 1204, 4, 128'h40300000000000000000000d546);
sram_add_entry(0, 6, 1208, 4, 128'h4030000000000000000000068ce);
sram_add_entry(0, 6, 1212, 4, 128'h40300000000000000000000ec8a);
sram_add_entry(0, 6, 1216, 4, 128'h40300000000000000000000fb29);
sram_add_entry(0, 6, 1220, 4, 128'h403000000000000000000000c7a);
sram_add_entry(0, 6, 1224, 4, 128'h403000000000000000000004760);
sram_add_entry(0, 6, 1228, 4, 128'h4030000000000000000000034fc);
sram_add_entry(0, 6, 1232, 4, 128'h403000000000000000000007313);
sram_add_entry(0, 6, 1236, 4, 128'h40300000000000000000000a699);
sram_add_entry(0, 6, 1240, 4, 128'h40300000000000000000000d724);
sram_add_entry(0, 6, 1244, 4, 128'h40300000000000000000000d427);
sram_add_entry(0, 6, 1248, 4, 128'h40300000000000000000000efcd);
sram_add_entry(0, 6, 1252, 4, 128'h40300000000000000000000f203);
sram_add_entry(0, 6, 1256, 4, 128'h4030000000000000000000041da);
sram_add_entry(0, 6, 1260, 4, 128'h40300000000000000000000390c);
sram_add_entry(0, 6, 1264, 4, 128'h403000000000000000000004b5a);
sram_add_entry(0, 6, 1268, 4, 128'h40300000000000000000000c980);
sram_add_entry(0, 6, 1272, 4, 128'h40300000000000000000000f62d);
sram_add_entry(0, 6, 1276, 4, 128'h403000000000000000000006fe6);
sram_add_entry(0, 6, 1280, 4, 128'h403000000000000000000008e36);
sram_add_entry(0, 6, 1284, 4, 128'h4030000000000000000000032cc);
sram_add_entry(0, 6, 1288, 4, 128'h40300000000000000000000ab0e);
sram_add_entry(0, 6, 1292, 4, 128'h4030000000000000000000087e8);
sram_add_entry(0, 6, 1296, 4, 128'h40300000000000000000000c504);
sram_add_entry(0, 6, 1300, 4, 128'h403000000000000000000002a99);
sram_add_entry(0, 6, 1304, 4, 128'h403000000000000000000006e23);
sram_add_entry(0, 6, 1308, 4, 128'h403000000000000000000007936);
sram_add_entry(0, 6, 1312, 4, 128'h40300000000000000000000e3be);
sram_add_entry(0, 6, 1316, 4, 128'h403000000000000000000003d8c);
sram_add_entry(0, 6, 1320, 4, 128'h40300000000000000000000689f);
sram_add_entry(0, 6, 1324, 4, 128'h40300000000000000000000d3c9);
sram_add_entry(0, 6, 1328, 4, 128'h40300000000000000000000cf80);
sram_add_entry(0, 6, 1332, 4, 128'h40300000000000000000000c8b4);
sram_add_entry(0, 6, 1336, 4, 128'h403000000000000000000007438);
sram_add_entry(0, 6, 1340, 4, 128'h40300000000000000000000d02d);
sram_add_entry(0, 6, 1344, 4, 128'h403000000000000000000005653);
sram_add_entry(0, 6, 1348, 4, 128'h40300000000000000000000462a);
sram_add_entry(0, 6, 1352, 4, 128'h4030000000000000000000079b6);
sram_add_entry(0, 6, 1356, 4, 128'h40300000000000000000000ff26);
sram_add_entry(0, 6, 1360, 4, 128'h40300000000000000000000c9f8);
sram_add_entry(0, 6, 1364, 4, 128'h40300000000000000000000c4de);
sram_add_entry(0, 6, 1368, 4, 128'h40300000000000000000000fd4b);
sram_add_entry(0, 6, 1372, 4, 128'h403000000000000000000001cc0);
sram_add_entry(0, 6, 1376, 4, 128'h403000000000000000000003961);
sram_add_entry(0, 6, 1380, 4, 128'h40300000000000000000000fac3);
sram_add_entry(0, 6, 1384, 4, 128'h4030000000000000000000096b3);
sram_add_entry(0, 6, 1388, 4, 128'h403000000000000000000001d75);
sram_add_entry(0, 6, 1392, 4, 128'h40300000000000000000000feeb);
sram_add_entry(0, 6, 1396, 4, 128'h403000000000000000000000d35);
sram_add_entry(0, 6, 1400, 4, 128'h40300000000000000000000c987);
sram_add_entry(0, 6, 1404, 4, 128'h403000000000000000000003659);
sram_add_entry(0, 6, 1408, 4, 128'h40300000000000000000000ed9a);
sram_add_entry(0, 6, 1412, 4, 128'h40300000000000000000000a77d);
sram_add_entry(0, 6, 1416, 4, 128'h4030000000000000000000000ea);
sram_add_entry(0, 6, 1420, 4, 128'h403000000000000000000006d0c);
sram_add_entry(0, 6, 1424, 4, 128'h403000000000000000000005f79);
sram_add_entry(0, 6, 1428, 4, 128'h403000000000000000000003ab0);
sram_add_entry(0, 6, 1432, 4, 128'h40300000000000000000000977e);
sram_add_entry(0, 6, 1436, 4, 128'h403000000000000000000003413);
sram_add_entry(0, 6, 1440, 4, 128'h40300000000000000000000990c);
sram_add_entry(0, 6, 1444, 4, 128'h40300000000000000000000530f);
sram_add_entry(0, 6, 1448, 4, 128'h403000000000000000000009949);
sram_add_entry(0, 6, 1452, 4, 128'h40300000000000000000000e132);
sram_add_entry(0, 6, 1456, 4, 128'h4030000000000000000000047e1);
sram_add_entry(0, 6, 1460, 4, 128'h4030000000000000000000077a2);
sram_add_entry(0, 6, 1464, 4, 128'h40300000000000000000000b608);
sram_add_entry(0, 6, 1468, 4, 128'h40300000000000000000000a7e7);
sram_add_entry(0, 6, 1472, 4, 128'h40300000000000000000000d940);
sram_add_entry(0, 6, 1476, 4, 128'h40300000000000000000000fb69);
sram_add_entry(0, 6, 1480, 4, 128'h40300000000000000000000131c);
sram_add_entry(0, 6, 1484, 4, 128'h403000000000000000000005d26);
sram_add_entry(0, 6, 1488, 4, 128'h40300000000000000000000a9cc);
sram_add_entry(0, 6, 1492, 4, 128'h403000000000000000000003677);
sram_add_entry(0, 6, 1496, 4, 128'h403000000000000000000004a66);
sram_add_entry(0, 6, 1500, 4, 128'h403000000000000000000009b09);
sram_add_entry(0, 6, 1504, 4, 128'h403000000000000000000003cea);
sram_add_entry(0, 6, 1508, 4, 128'h403000000000000000000004f86);
sram_add_entry(0, 6, 1512, 4, 128'h403000000000000000000005443);
sram_add_entry(0, 6, 1516, 4, 128'h40300000000000000000000cc10);
sram_add_entry(0, 6, 1520, 4, 128'h40300000000000000000000a83c);
sram_add_entry(0, 6, 1524, 4, 128'h403000000000000000000002399);
sram_add_entry(0, 6, 1528, 4, 128'h40300000000000000000000eed1);
sram_add_entry(0, 6, 1532, 4, 128'h403000000000000000000008b00);
sram_add_entry(0, 6, 1536, 4, 128'h40300000000000000000000c875);
sram_add_entry(0, 6, 1540, 4, 128'h4030000000000000000000030e5);
sram_add_entry(0, 6, 1544, 4, 128'h40300000000000000000000c912);
sram_add_entry(0, 6, 1548, 4, 128'h4030000000000000000000095c2);
sram_add_entry(0, 6, 1552, 4, 128'h40300000000000000000000f263);
sram_add_entry(0, 6, 1556, 4, 128'h403000000000000000000005500);
sram_add_entry(0, 6, 1560, 4, 128'h403000000000000000000003863);
sram_add_entry(0, 6, 1564, 4, 128'h40300000000000000000000da52);
sram_add_entry(0, 6, 1568, 4, 128'h403000000000000000000004a7f);
sram_add_entry(0, 6, 1572, 4, 128'h40300000000000000000000031b);
sram_add_entry(0, 6, 1576, 4, 128'h403000000000000000000001bac);
sram_add_entry(0, 6, 1580, 4, 128'h403000000000000000000009b43);
sram_add_entry(0, 6, 1584, 4, 128'h40300000000000000000000a30f);
sram_add_entry(0, 6, 1588, 4, 128'h40300000000000000000000c88d);
sram_add_entry(0, 6, 1592, 4, 128'h403000000000000000000001146);
sram_add_entry(0, 6, 1596, 4, 128'h4030000000000000000000033e3);
sram_add_entry(0, 6, 1600, 4, 128'h40300000000000000000000d222);
sram_add_entry(0, 6, 1604, 4, 128'h40300000000000000000000bf0a);
sram_add_entry(0, 6, 1608, 4, 128'h403000000000000000000008d89);
sram_add_entry(0, 6, 1612, 4, 128'h4030000000000000000000024f0);
sram_add_entry(0, 6, 1616, 4, 128'h403000000000000000000000e2e);
sram_add_entry(0, 6, 1620, 4, 128'h40300000000000000000000d40c);
sram_add_entry(0, 6, 1624, 4, 128'h403000000000000000000002570);
sram_add_entry(0, 6, 1628, 4, 128'h403000000000000000000002acc);
sram_add_entry(0, 6, 1632, 4, 128'h403000000000000000000003dc1);
sram_add_entry(0, 6, 1636, 4, 128'h403000000000000000000005b5b);
sram_add_entry(0, 6, 1640, 4, 128'h403000000000000000000004198);
sram_add_entry(0, 6, 1644, 4, 128'h403000000000000000000008e6d);
sram_add_entry(0, 6, 1648, 4, 128'h4030000000000000000000012a8);
sram_add_entry(0, 6, 1652, 4, 128'h40300000000000000000000fd89);
sram_add_entry(0, 6, 1656, 4, 128'h403000000000000000000002577);
sram_add_entry(0, 6, 1660, 4, 128'h403000000000000000000003edf);
sram_add_entry(0, 6, 1664, 4, 128'h403000000000000000000006331);
sram_add_entry(0, 6, 1668, 4, 128'h403000000000000000000004747);
sram_add_entry(0, 6, 1672, 4, 128'h403000000000000000000002327);
sram_add_entry(0, 6, 1676, 4, 128'h403000000000000000000004c09);
sram_add_entry(0, 6, 1680, 4, 128'h403000000000000000000001a17);
sram_add_entry(0, 6, 1684, 4, 128'h40300000000000000000000a395);
sram_add_entry(0, 6, 1688, 4, 128'h403000000000000000000000c94);
sram_add_entry(0, 6, 1692, 4, 128'h403000000000000000000000174);
sram_add_entry(0, 6, 1696, 4, 128'h40300000000000000000000212e);
sram_add_entry(0, 6, 1700, 4, 128'h4030000000000000000000080ab);
sram_add_entry(0, 6, 1704, 4, 128'h40300000000000000000000a361);
sram_add_entry(0, 6, 1708, 4, 128'h40300000000000000000000fbf6);
sram_add_entry(0, 6, 1712, 4, 128'h40300000000000000000000d291);
sram_add_entry(0, 6, 1716, 4, 128'h4030000000000000000000081bf);
sram_add_entry(0, 6, 1720, 4, 128'h403000000000000000000000c9e);
sram_add_entry(0, 6, 1724, 4, 128'h40300000000000000000000e846);
sram_add_entry(0, 6, 1728, 4, 128'h403000000000000000000000d5c);
sram_add_entry(0, 6, 1732, 4, 128'h40300000000000000000000ce2a);
sram_add_entry(0, 6, 1736, 4, 128'h40300000000000000000000fa53);
sram_add_entry(0, 6, 1740, 4, 128'h403000000000000000000004afe);
sram_add_entry(0, 6, 1744, 4, 128'h40300000000000000000000215d);
sram_add_entry(0, 6, 1748, 4, 128'h40300000000000000000000a8f9);
sram_add_entry(0, 6, 1752, 4, 128'h403000000000000000000009fff);
sram_add_entry(0, 6, 1756, 4, 128'h40300000000000000000000539d);
sram_add_entry(0, 6, 1760, 4, 128'h403000000000000000000002c1e);
sram_add_entry(0, 6, 1764, 4, 128'h403000000000000000000003ea8);
sram_add_entry(0, 6, 1768, 4, 128'h403000000000000000000008d4c);
sram_add_entry(0, 6, 1772, 4, 128'h403000000000000000000009c5c);
sram_add_entry(0, 6, 1776, 4, 128'h40300000000000000000000db37);
sram_add_entry(0, 6, 1780, 4, 128'h40300000000000000000000a769);
sram_add_entry(0, 6, 1784, 4, 128'h403000000000000000000001c12);
sram_add_entry(0, 6, 1788, 4, 128'h4030000000000000000000042e3);
sram_add_entry(0, 6, 1792, 4, 128'h40300000000000000000000c8ca);
sram_add_entry(0, 6, 1796, 4, 128'h40300000000000000000000acf8);
sram_add_entry(0, 6, 1800, 4, 128'h40300000000000000000000f770);
sram_add_entry(0, 6, 1804, 4, 128'h4030000000000000000000057ff);
sram_add_entry(0, 6, 1808, 4, 128'h403000000000000000000006a40);
sram_add_entry(0, 6, 1812, 4, 128'h403000000000000000000006579);
sram_add_entry(0, 6, 1816, 4, 128'h40300000000000000000000499e);
sram_add_entry(0, 6, 1820, 4, 128'h4030000000000000000000027a1);
sram_add_entry(0, 6, 1824, 4, 128'h403000000000000000000009123);
sram_add_entry(0, 6, 1828, 4, 128'h40300000000000000000000a641);
sram_add_entry(0, 6, 1832, 4, 128'h4030000000000000000000080db);
sram_add_entry(0, 6, 1836, 4, 128'h40300000000000000000000cbf3);
sram_add_entry(0, 6, 1840, 4, 128'h40300000000000000000000a9a5);
sram_add_entry(0, 6, 1844, 4, 128'h403000000000000000000003824);
sram_add_entry(0, 6, 1848, 4, 128'h40300000000000000000000c25d);
sram_add_entry(0, 6, 1852, 4, 128'h40300000000000000000000d240);
sram_add_entry(0, 6, 1856, 4, 128'h40300000000000000000000bebd);
sram_add_entry(0, 6, 1860, 4, 128'h40300000000000000000000e5fc);
sram_add_entry(0, 6, 1864, 4, 128'h403000000000000000000007e08);
sram_add_entry(0, 6, 1868, 4, 128'h403000000000000000000006999);
sram_add_entry(0, 6, 1872, 4, 128'h40300000000000000000000a30b);
sram_add_entry(0, 6, 1876, 4, 128'h40300000000000000000000b086);
sram_add_entry(0, 6, 1880, 4, 128'h403000000000000000000002c3e);
sram_add_entry(0, 6, 1884, 4, 128'h40300000000000000000000e232);
sram_add_entry(0, 6, 1888, 4, 128'h40300000000000000000000c378);
sram_add_entry(0, 6, 1892, 4, 128'h40300000000000000000000b14c);
sram_add_entry(0, 6, 1896, 4, 128'h403000000000000000000002bb7);
sram_add_entry(0, 6, 1900, 4, 128'h403000000000000000000000d28);
sram_add_entry(0, 6, 1904, 4, 128'h40300000000000000000000b678);
sram_add_entry(0, 6, 1908, 4, 128'h40300000000000000000000a845);
sram_add_entry(0, 6, 1912, 4, 128'h40300000000000000000000c805);
sram_add_entry(0, 6, 1916, 4, 128'h40300000000000000000000f905);
sram_add_entry(0, 6, 1920, 4, 128'h403000000000000000000005909);
sram_add_entry(0, 6, 1924, 4, 128'h403000000000000000000001850);
sram_add_entry(0, 6, 1928, 4, 128'h403000000000000000000003708);
sram_add_entry(0, 6, 1932, 4, 128'h403000000000000000000003bb1);
sram_add_entry(0, 6, 1936, 4, 128'h40300000000000000000000fe35);
sram_add_entry(0, 6, 1940, 4, 128'h403000000000000000000003010);
sram_add_entry(0, 6, 1944, 4, 128'h40300000000000000000000222f);
sram_add_entry(0, 6, 1948, 4, 128'h4030000000000000000000056fa);
sram_add_entry(0, 6, 1952, 4, 128'h403000000000000000000003023);
sram_add_entry(0, 6, 1956, 4, 128'h40300000000000000000000de51);
sram_add_entry(0, 6, 1960, 4, 128'h403000000000000000000009900);
sram_add_entry(0, 6, 1964, 4, 128'h403000000000000000000007b27);
sram_add_entry(0, 6, 1968, 4, 128'h40300000000000000000000a678);
sram_add_entry(0, 6, 1972, 4, 128'h403000000000000000000004ff3);
sram_add_entry(0, 6, 1976, 4, 128'h4030000000000000000000095fc);
sram_add_entry(0, 6, 1980, 4, 128'h403000000000000000000008d2c);
sram_add_entry(0, 6, 1984, 4, 128'h403000000000000000000008a9e);
sram_add_entry(0, 6, 1988, 4, 128'h403000000000000000000000eef);
sram_add_entry(0, 6, 1992, 4, 128'h40300000000000000000000d8e7);
sram_add_entry(0, 6, 1996, 4, 128'h403000000000000000000000a7e);
sram_add_entry(0, 6, 2000, 4, 128'h4030000000000000000000019a1);
sram_add_entry(0, 6, 2004, 4, 128'h40300000000000000000000ec33);
sram_add_entry(0, 6, 2008, 4, 128'h40300000000000000000000a05a);
sram_add_entry(0, 6, 2012, 4, 128'h403000000000000000000007046);
sram_add_entry(0, 6, 2016, 4, 128'h403000000000000000000002ea1);
sram_add_entry(0, 6, 2020, 4, 128'h403000000000000000000009bf1);
sram_add_entry(0, 6, 2024, 4, 128'h40300000000000000000000ac89);
sram_add_entry(0, 6, 2028, 4, 128'h403000000000000000000001572);
sram_add_entry(0, 6, 2032, 4, 128'h403000000000000000000001b4c);
sram_add_entry(0, 6, 2036, 4, 128'h4030000000000000000000066b0);
sram_add_entry(0, 6, 2040, 4, 128'h40300000000000000000000046e);
sram_add_entry(0, 6, 2044, 4, 128'h40300000000000000000000f521);
sram_add_entry(0, 6, 2048, 4, 128'h403000000000000000000007fed);
sram_add_entry(0, 6, 2052, 4, 128'h40300000000000000000000a538);
sram_add_entry(0, 6, 2056, 4, 128'h40300000000000000000000721d);
sram_add_entry(0, 6, 2060, 4, 128'h403000000000000000000001f85);
sram_add_entry(0, 6, 2064, 4, 128'h40300000000000000000000ddcf);
sram_add_entry(0, 6, 2068, 4, 128'h40300000000000000000000923c);
sram_add_entry(0, 6, 2072, 4, 128'h403000000000000000000005be3);
sram_add_entry(0, 6, 2076, 4, 128'h40300000000000000000000c41c);
sram_add_entry(0, 6, 2080, 4, 128'h403000000000000000000000e73);
sram_add_entry(0, 6, 2084, 4, 128'h403000000000000000000004046);
sram_add_entry(0, 6, 2088, 4, 128'h403000000000000000000008109);
sram_add_entry(0, 6, 2092, 4, 128'h40300000000000000000000966e);
sram_add_entry(0, 6, 2096, 4, 128'h40300000000000000000000e61a);
sram_add_entry(0, 6, 2100, 4, 128'h403000000000000000000007975);
sram_add_entry(0, 6, 2104, 4, 128'h40300000000000000000000d88c);
sram_add_entry(0, 6, 2108, 4, 128'h40300000000000000000000645a);
sram_add_entry(0, 6, 2112, 4, 128'h4030000000000000000000087d2);
sram_add_entry(0, 6, 2116, 4, 128'h40300000000000000000000619d);
sram_add_entry(0, 6, 2120, 4, 128'h4030000000000000000000093fc);
sram_add_entry(0, 6, 2124, 4, 128'h403000000000000000000001d1b);
sram_add_entry(0, 6, 2128, 4, 128'h40300000000000000000000e191);
sram_add_entry(0, 6, 2132, 4, 128'h403000000000000000000008160);
sram_add_entry(0, 6, 2136, 4, 128'h40300000000000000000000fd5e);
sram_add_entry(0, 6, 2140, 4, 128'h40300000000000000000000ad9e);
sram_add_entry(0, 6, 2144, 4, 128'h40300000000000000000000e6bc);
sram_add_entry(0, 6, 2148, 4, 128'h403000000000000000000009199);
sram_add_entry(0, 6, 2152, 4, 128'h40300000000000000000000ffde);
sram_add_entry(0, 6, 2156, 4, 128'h403000000000000000000006c77);
sram_add_entry(0, 6, 2160, 4, 128'h403000000000000000000004d6c);
sram_add_entry(0, 6, 2164, 4, 128'h40300000000000000000000d10a);
sram_add_entry(0, 6, 2168, 4, 128'h40300000000000000000000e977);
sram_add_entry(0, 6, 2172, 4, 128'h403000000000000000000004135);
sram_add_entry(0, 6, 2176, 4, 128'h40300000000000000000000bcb9);
sram_add_entry(0, 6, 2180, 4, 128'h40300000000000000000000a3ed);
sram_add_entry(0, 6, 2184, 4, 128'h4030000000000000000000081ec);
sram_add_entry(0, 6, 2188, 4, 128'h4030000000000000000000040f1);
sram_add_entry(0, 6, 2192, 4, 128'h40300000000000000000000e12e);
sram_add_entry(0, 6, 2196, 4, 128'h403000000000000000000008bd3);
sram_add_entry(0, 6, 2200, 4, 128'h4030000000000000000000005de);
sram_add_entry(0, 6, 2204, 4, 128'h40300000000000000000000852e);
sram_add_entry(0, 6, 2208, 4, 128'h4030000000000000000000089be);
sram_add_entry(0, 6, 2212, 4, 128'h403000000000000000000009c0c);
sram_add_entry(0, 6, 2216, 4, 128'h4030000000000000000000058fb);
sram_add_entry(0, 6, 2220, 4, 128'h40300000000000000000000aa88);
sram_add_entry(0, 6, 2224, 4, 128'h40300000000000000000000b6f4);
sram_add_entry(0, 6, 2228, 4, 128'h403000000000000000000005206);
sram_add_entry(0, 6, 2232, 4, 128'h403000000000000000000006efd);
sram_add_entry(0, 6, 2236, 4, 128'h40300000000000000000000432b);
sram_add_entry(0, 6, 2240, 4, 128'h40300000000000000000000715e);
sram_add_entry(0, 6, 2244, 4, 128'h403000000000000000000000633);
sram_add_entry(0, 6, 2248, 4, 128'h403000000000000000000009f03);
sram_add_entry(0, 6, 2252, 4, 128'h40300000000000000000000ed63);
sram_add_entry(0, 6, 2256, 4, 128'h403000000000000000000007a86);
sram_add_entry(0, 6, 2260, 4, 128'h403000000000000000000008df8);
sram_add_entry(0, 6, 2264, 4, 128'h403000000000000000000004007);
sram_add_entry(0, 6, 2268, 4, 128'h40300000000000000000000db34);
sram_add_entry(0, 6, 2272, 4, 128'h403000000000000000000007aa9);
sram_add_entry(0, 6, 2276, 4, 128'h4030000000000000000000074d0);
sram_add_entry(0, 6, 2280, 4, 128'h40300000000000000000000c8a5);
sram_add_entry(0, 6, 2284, 4, 128'h403000000000000000000002c9d);
sram_add_entry(0, 6, 2288, 4, 128'h403000000000000000000007b79);
sram_add_entry(0, 6, 2292, 4, 128'h40300000000000000000000f1d6);
sram_add_entry(0, 6, 2296, 4, 128'h403000000000000000000008452);
sram_add_entry(0, 6, 2300, 4, 128'h40300000000000000000000a758);
sram_add_entry(0, 6, 2304, 4, 128'h40300000000000000000000c377);
sram_add_entry(0, 6, 2308, 4, 128'h403000000000000000000009a0a);
sram_add_entry(0, 6, 2312, 4, 128'h4030000000000000000000051a0);
sram_add_entry(0, 6, 2316, 4, 128'h40300000000000000000000e2f5);
sram_add_entry(0, 6, 2320, 4, 128'h40300000000000000000000ebd0);
sram_add_entry(0, 6, 2324, 4, 128'h403000000000000000000000bba);
sram_add_entry(0, 6, 2328, 4, 128'h40300000000000000000000495a);
sram_add_entry(0, 6, 2332, 4, 128'h4030000000000000000000084ac);
sram_add_entry(0, 6, 2336, 4, 128'h403000000000000000000000d77);
sram_add_entry(0, 6, 2340, 4, 128'h40300000000000000000000ceef);
sram_add_entry(0, 6, 2344, 4, 128'h40300000000000000000000bb05);
sram_add_entry(0, 6, 2348, 4, 128'h403000000000000000000007e66);
sram_add_entry(0, 6, 2352, 4, 128'h403000000000000000000006e53);
sram_add_entry(0, 6, 2356, 4, 128'h403000000000000000000009083);
sram_add_entry(0, 6, 2360, 4, 128'h4030000000000000000000048cc);
sram_add_entry(0, 6, 2364, 4, 128'h403000000000000000000008be5);
sram_add_entry(0, 6, 2368, 4, 128'h403000000000000000000005f88);
sram_add_entry(0, 6, 2372, 4, 128'h4030000000000000000000068a8);
sram_add_entry(0, 6, 2376, 4, 128'h40300000000000000000000c805);
sram_add_entry(0, 6, 2380, 4, 128'h403000000000000000000009ecf);
sram_add_entry(0, 6, 2384, 4, 128'h40300000000000000000000d5f0);
sram_add_entry(0, 6, 2388, 4, 128'h403000000000000000000001cfc);
sram_add_entry(0, 6, 2392, 4, 128'h40300000000000000000000c265);
sram_add_entry(0, 6, 2396, 4, 128'h40300000000000000000000d9b4);
sram_add_entry(0, 6, 2400, 4, 128'h403000000000000000000005053);
sram_add_entry(0, 6, 2404, 4, 128'h403000000000000000000006860);
sram_add_entry(0, 6, 2408, 4, 128'h40300000000000000000000039a);
sram_add_entry(0, 6, 2412, 4, 128'h40300000000000000000000bb6c);
sram_add_entry(0, 6, 2416, 4, 128'h40300000000000000000000210c);
sram_add_entry(0, 6, 2420, 4, 128'h403000000000000000000006980);
sram_add_entry(0, 6, 2424, 4, 128'h40300000000000000000000a25d);
sram_add_entry(0, 6, 2428, 4, 128'h403000000000000000000009aec);
sram_add_entry(0, 6, 2432, 4, 128'h40300000000000000000000b8c5);
sram_add_entry(0, 6, 2436, 4, 128'h40300000000000000000000a45b);
sram_add_entry(0, 6, 2440, 4, 128'h403000000000000000000001bfb);
sram_add_entry(0, 6, 2444, 4, 128'h4030000000000000000000058d3);
sram_add_entry(0, 6, 2448, 4, 128'h403000000000000000000000e69);
sram_add_entry(0, 6, 2452, 4, 128'h403000000000000000000002820);
sram_add_entry(0, 6, 2456, 4, 128'h403000000000000000000004054);
sram_add_entry(0, 6, 2460, 4, 128'h40300000000000000000000b2e2);
sram_add_entry(0, 6, 2464, 4, 128'h403000000000000000000000316);
sram_add_entry(0, 6, 2468, 4, 128'h403000000000000000000007aa9);
sram_add_entry(0, 6, 2472, 4, 128'h4030000000000000000000010a8);
sram_add_entry(0, 6, 2476, 4, 128'h40300000000000000000000e18a);
sram_add_entry(0, 6, 2480, 4, 128'h40300000000000000000000ab13);
sram_add_entry(0, 6, 2484, 4, 128'h40300000000000000000000f1d1);
sram_add_entry(0, 6, 2488, 4, 128'h4030000000000000000000014f2);
sram_add_entry(0, 6, 2492, 4, 128'h403000000000000000000006822);
sram_add_entry(0, 6, 2496, 4, 128'h403000000000000000000004228);
sram_add_entry(0, 6, 2500, 4, 128'h4030000000000000000000081e5);
sram_add_entry(0, 6, 2504, 4, 128'h403000000000000000000006203);
sram_add_entry(0, 6, 2508, 4, 128'h4030000000000000000000048b2);
sram_add_entry(0, 6, 2512, 4, 128'h403000000000000000000007b40);
sram_add_entry(0, 6, 2516, 4, 128'h40300000000000000000000f692);
sram_add_entry(0, 6, 2520, 4, 128'h40300000000000000000000ab7e);
sram_add_entry(0, 6, 2524, 4, 128'h40300000000000000000000ce0c);
sram_add_entry(0, 6, 2528, 4, 128'h40300000000000000000000a40b);
sram_add_entry(0, 6, 2532, 4, 128'h403000000000000000000004636);
sram_add_entry(0, 6, 2536, 4, 128'h403000000000000000000003aee);
sram_add_entry(0, 6, 2540, 4, 128'h40300000000000000000000ef6c);
sram_add_entry(0, 6, 2544, 4, 128'h40300000000000000000000928f);
sram_add_entry(0, 6, 2548, 4, 128'h40300000000000000000000d60f);
sram_add_entry(0, 6, 2552, 4, 128'h40300000000000000000000bd68);
sram_add_entry(0, 6, 2556, 4, 128'h4030000000000000000000030c9);
sram_add_entry(0, 6, 2560, 4, 128'h40300000000000000000000cbd2);
sram_add_entry(0, 6, 2564, 4, 128'h40300000000000000000000d53c);
sram_add_entry(0, 6, 2568, 4, 128'h403000000000000000000001685);
sram_add_entry(0, 6, 2572, 4, 128'h403000000000000000000002195);
sram_add_entry(0, 6, 2576, 4, 128'h40300000000000000000000a4e0);
sram_add_entry(0, 6, 2580, 4, 128'h40300000000000000000000aede);
sram_add_entry(0, 6, 2584, 4, 128'h40300000000000000000000b476);
sram_add_entry(0, 6, 2588, 4, 128'h403000000000000000000004bdf);
sram_add_entry(0, 6, 2592, 4, 128'h403000000000000000000003cb8);
sram_add_entry(0, 6, 2596, 4, 128'h40300000000000000000000d010);
sram_add_entry(0, 6, 2600, 4, 128'h40300000000000000000000946b);
sram_add_entry(0, 6, 2604, 4, 128'h40300000000000000000000afd1);
sram_add_entry(0, 6, 2608, 4, 128'h40300000000000000000000f204);
sram_add_entry(0, 6, 2612, 4, 128'h403000000000000000000006781);
sram_add_entry(0, 6, 2616, 4, 128'h40300000000000000000000b5f3);
sram_add_entry(0, 6, 2620, 4, 128'h40300000000000000000000a278);
sram_add_entry(0, 6, 2624, 4, 128'h403000000000000000000004a51);
sram_add_entry(0, 6, 2628, 4, 128'h40300000000000000000000f899);
sram_add_entry(0, 6, 2632, 4, 128'h40300000000000000000000ed90);
sram_add_entry(0, 6, 2636, 4, 128'h40300000000000000000000edf8);
sram_add_entry(0, 6, 2640, 4, 128'h40300000000000000000000252e);
sram_add_entry(0, 6, 2644, 4, 128'h4030000000000000000000052aa);
sram_add_entry(0, 6, 2648, 4, 128'h40300000000000000000000162b);
sram_add_entry(0, 6, 2652, 4, 128'h40300000000000000000000fbd9);
sram_add_entry(0, 6, 2656, 4, 128'h4030000000000000000000012df);
sram_add_entry(0, 6, 2660, 4, 128'h403000000000000000000007022);
sram_add_entry(0, 6, 2664, 4, 128'h403000000000000000000001a1f);
sram_add_entry(0, 6, 2668, 4, 128'h40300000000000000000000f03f);
sram_add_entry(0, 6, 2672, 4, 128'h403000000000000000000000324);
sram_add_entry(0, 6, 2676, 4, 128'h40300000000000000000000962c);
sram_add_entry(0, 6, 2680, 4, 128'h403000000000000000000003723);
sram_add_entry(0, 6, 2684, 4, 128'h403000000000000000000007c70);
sram_add_entry(0, 6, 2688, 4, 128'h403000000000000000000004bc5);
sram_add_entry(0, 6, 2692, 4, 128'h40300000000000000000000ca6b);
sram_add_entry(0, 6, 2696, 4, 128'h403000000000000000000006f8b);
sram_add_entry(0, 6, 2700, 4, 128'h403000000000000000000004565);
sram_add_entry(0, 6, 2704, 4, 128'h403000000000000000000003366);
sram_add_entry(0, 6, 2708, 4, 128'h40300000000000000000000e66a);
sram_add_entry(0, 6, 2712, 4, 128'h403000000000000000000000209);
sram_add_entry(0, 6, 2716, 4, 128'h40300000000000000000000c785);
sram_add_entry(0, 6, 2720, 4, 128'h40300000000000000000000dff4);
sram_add_entry(0, 6, 2724, 4, 128'h40300000000000000000000050e);
sram_add_entry(0, 6, 2728, 4, 128'h40300000000000000000000a9f5);
sram_add_entry(0, 6, 2732, 4, 128'h40300000000000000000000ba20);
sram_add_entry(0, 6, 2736, 4, 128'h40300000000000000000000ba1d);
sram_add_entry(0, 6, 2740, 4, 128'h40300000000000000000000a04d);
sram_add_entry(0, 6, 2744, 4, 128'h403000000000000000000005474);
sram_add_entry(0, 6, 2748, 4, 128'h403000000000000000000004961);
sram_add_entry(0, 6, 2752, 4, 128'h40300000000000000000000b74e);
sram_add_entry(0, 6, 2756, 4, 128'h40300000000000000000000e69a);
sram_add_entry(0, 6, 2760, 4, 128'h40300000000000000000000e108);
sram_add_entry(0, 6, 2764, 4, 128'h4030000000000000000000088aa);
sram_add_entry(0, 6, 2768, 4, 128'h40300000000000000000000d5b3);
sram_add_entry(0, 6, 2772, 4, 128'h40300000000000000000000bb4c);
sram_add_entry(0, 6, 2776, 4, 128'h403000000000000000000009ba6);
sram_add_entry(0, 6, 2780, 4, 128'h403000000000000000000004930);
sram_add_entry(0, 6, 2784, 4, 128'h40300000000000000000000e153);
sram_add_entry(0, 6, 2788, 4, 128'h403000000000000000000002cbf);
sram_add_entry(0, 6, 2792, 4, 128'h40300000000000000000000f52a);
sram_add_entry(0, 6, 2796, 4, 128'h40300000000000000000000e6da);
sram_add_entry(0, 6, 2800, 4, 128'h40300000000000000000000e180);
sram_add_entry(0, 2, 0, 4, 128'h7ab000000000000000000deadbf);
sram_add_entry(0, 2, 4, 4, 128'h40300000000000000000000c153);
sram_add_entry(0, 2, 8, 4, 128'h40300000000000000000000df3d);
sram_add_entry(0, 2, 12, 4, 128'h403000000000000000000003f56);
sram_add_entry(0, 2, 16, 4, 128'h40300000000000000000000b758);
sram_add_entry(0, 2, 20, 4, 128'h40300000000000000000000972b);
sram_add_entry(0, 2, 24, 4, 128'h40300000000000000000000624e);
sram_add_entry(0, 2, 28, 4, 128'h40300000000000000000000d51d);
sram_add_entry(0, 2, 32, 4, 128'h40300000000000000000000b905);
sram_add_entry(0, 2, 36, 4, 128'h40300000000000000000000a8a9);
sram_add_entry(0, 2, 40, 4, 128'h40300000000000000000000a7c9);
sram_add_entry(0, 2, 44, 4, 128'h4030000000000000000000037f8);
sram_add_entry(0, 2, 48, 4, 128'h40300000000000000000000ee8c);
sram_add_entry(0, 2, 52, 4, 128'h4030000000000000000000095f5);
sram_add_entry(0, 2, 56, 4, 128'h40300000000000000000000be40);
sram_add_entry(0, 2, 60, 4, 128'h40300000000000000000000a2c3);
sram_add_entry(0, 2, 64, 4, 128'h403000000000000000000003275);
sram_add_entry(0, 2, 68, 4, 128'h40300000000000000000000f5ff);
sram_add_entry(0, 2, 72, 4, 128'h4030000000000000000000084c6);
sram_add_entry(0, 2, 76, 4, 128'h40300000000000000000000a54c);
sram_add_entry(0, 2, 80, 4, 128'h40300000000000000000000c4f3);
sram_add_entry(0, 2, 84, 4, 128'h403000000000000000000004a8d);
sram_add_entry(0, 2, 88, 4, 128'h40300000000000000000000fe35);
sram_add_entry(0, 2, 92, 4, 128'h40300000000000000000000dff6);
sram_add_entry(0, 2, 96, 4, 128'h403000000000000000000001765);
sram_add_entry(0, 2, 100, 4, 128'h40300000000000000000000b292);
sram_add_entry(0, 2, 104, 4, 128'h403000000000000000000004d71);
sram_add_entry(0, 2, 108, 4, 128'h403000000000000000000004d83);
sram_add_entry(0, 2, 112, 4, 128'h403000000000000000000006c69);
sram_add_entry(0, 2, 116, 4, 128'h403000000000000000000001c6b);
sram_add_entry(0, 2, 120, 4, 128'h40300000000000000000000a4bb);
sram_add_entry(0, 2, 124, 4, 128'h403000000000000000000009c42);
sram_add_entry(0, 2, 128, 4, 128'h40300000000000000000000f399);
sram_add_entry(0, 2, 132, 4, 128'h40300000000000000000000e276);
sram_add_entry(0, 2, 136, 4, 128'h40300000000000000000000782c);
sram_add_entry(0, 2, 140, 4, 128'h403000000000000000000000556);
sram_add_entry(0, 2, 144, 4, 128'h403000000000000000000003d19);
sram_add_entry(0, 2, 148, 4, 128'h4030000000000000000000061df);
sram_add_entry(0, 2, 152, 4, 128'h4030000000000000000000025c0);
sram_add_entry(0, 2, 156, 4, 128'h403000000000000000000004c4b);
sram_add_entry(0, 2, 160, 4, 128'h403000000000000000000000962);
sram_add_entry(0, 2, 164, 4, 128'h40300000000000000000000a4e4);
sram_add_entry(0, 2, 168, 4, 128'h403000000000000000000003376);
sram_add_entry(0, 2, 172, 4, 128'h40300000000000000000000bfd6);
sram_add_entry(0, 2, 176, 4, 128'h403000000000000000000002121);
sram_add_entry(0, 2, 180, 4, 128'h40300000000000000000000393a);
sram_add_entry(0, 2, 184, 4, 128'h40300000000000000000000c59c);
sram_add_entry(0, 2, 188, 4, 128'h40300000000000000000000bab5);
sram_add_entry(0, 2, 192, 4, 128'h403000000000000000000004d89);
sram_add_entry(0, 2, 196, 4, 128'h4030000000000000000000078ec);
sram_add_entry(0, 2, 200, 4, 128'h403000000000000000000009051);
sram_add_entry(0, 2, 204, 4, 128'h403000000000000000000001fb5);
sram_add_entry(0, 2, 208, 4, 128'h4030000000000000000000084c3);
sram_add_entry(0, 2, 212, 4, 128'h40300000000000000000000532f);
sram_add_entry(0, 2, 216, 4, 128'h40300000000000000000000fcec);
sram_add_entry(0, 2, 220, 4, 128'h40300000000000000000000460e);
sram_add_entry(0, 2, 224, 4, 128'h4030000000000000000000012a9);
sram_add_entry(0, 2, 228, 4, 128'h403000000000000000000002f22);
sram_add_entry(0, 2, 232, 4, 128'h40300000000000000000000297d);
sram_add_entry(0, 2, 236, 4, 128'h403000000000000000000002f95);
sram_add_entry(0, 2, 240, 4, 128'h403000000000000000000003952);
sram_add_entry(0, 2, 244, 4, 128'h4030000000000000000000059e5);
sram_add_entry(0, 2, 248, 4, 128'h403000000000000000000004201);
sram_add_entry(0, 2, 252, 4, 128'h40300000000000000000000abfb);
sram_add_entry(0, 2, 256, 4, 128'h40300000000000000000000890f);
sram_add_entry(0, 2, 260, 4, 128'h40300000000000000000000fc14);
sram_add_entry(0, 2, 264, 4, 128'h40300000000000000000000561d);
sram_add_entry(0, 2, 268, 4, 128'h403000000000000000000009b06);
sram_add_entry(0, 2, 272, 4, 128'h403000000000000000000000c82);
sram_add_entry(0, 2, 276, 4, 128'h403000000000000000000007392);
sram_add_entry(0, 2, 280, 4, 128'h4030000000000000000000069f8);
sram_add_entry(0, 2, 284, 4, 128'h40300000000000000000000ab52);
sram_add_entry(0, 2, 288, 4, 128'h4030000000000000000000046a7);
sram_add_entry(0, 2, 292, 4, 128'h4030000000000000000000088bd);
sram_add_entry(0, 2, 296, 4, 128'h40300000000000000000000b6c5);
sram_add_entry(0, 2, 300, 4, 128'h40300000000000000000000f611);
sram_add_entry(0, 2, 304, 4, 128'h403000000000000000000001778);
sram_add_entry(0, 2, 308, 4, 128'h403000000000000000000009317);
sram_add_entry(0, 2, 312, 4, 128'h40300000000000000000000b32f);
sram_add_entry(0, 2, 316, 4, 128'h40300000000000000000000f584);
sram_add_entry(0, 2, 320, 4, 128'h403000000000000000000001183);
sram_add_entry(0, 2, 324, 4, 128'h40300000000000000000000e56f);
sram_add_entry(0, 2, 328, 4, 128'h4030000000000000000000073f8);
sram_add_entry(0, 2, 332, 4, 128'h40300000000000000000000e077);
sram_add_entry(0, 2, 336, 4, 128'h403000000000000000000009ca6);
sram_add_entry(0, 2, 340, 4, 128'h403000000000000000000009acc);
sram_add_entry(0, 2, 344, 4, 128'h40300000000000000000000165c);
sram_add_entry(0, 2, 348, 4, 128'h40300000000000000000000956e);
sram_add_entry(0, 2, 352, 4, 128'h40300000000000000000000a541);
sram_add_entry(0, 2, 356, 4, 128'h40300000000000000000000b89e);
sram_add_entry(0, 2, 360, 4, 128'h403000000000000000000003001);
sram_add_entry(0, 2, 364, 4, 128'h4030000000000000000000023b7);
sram_add_entry(0, 2, 368, 4, 128'h40300000000000000000000a9b2);
sram_add_entry(0, 2, 372, 4, 128'h40300000000000000000000f128);
sram_add_entry(0, 2, 376, 4, 128'h40300000000000000000000b305);
sram_add_entry(0, 2, 380, 4, 128'h403000000000000000000000032);
sram_add_entry(0, 2, 384, 4, 128'h403000000000000000000001876);
sram_add_entry(0, 2, 388, 4, 128'h40300000000000000000000f881);
sram_add_entry(0, 2, 392, 4, 128'h40300000000000000000000dbfb);
sram_add_entry(0, 2, 396, 4, 128'h40300000000000000000000aa91);
sram_add_entry(0, 2, 400, 4, 128'h403000000000000000000004b52);
sram_add_entry(0, 2, 404, 4, 128'h40300000000000000000000b267);
sram_add_entry(0, 2, 408, 4, 128'h403000000000000000000007b38);
sram_add_entry(0, 2, 412, 4, 128'h403000000000000000000003af9);
sram_add_entry(0, 2, 416, 4, 128'h403000000000000000000001df7);
sram_add_entry(0, 2, 420, 4, 128'h40300000000000000000000f165);
sram_add_entry(0, 2, 424, 4, 128'h40300000000000000000000202f);
sram_add_entry(0, 2, 428, 4, 128'h4030000000000000000000040c4);
sram_add_entry(0, 2, 432, 4, 128'h403000000000000000000001275);
sram_add_entry(0, 2, 436, 4, 128'h4030000000000000000000067fe);
sram_add_entry(0, 2, 440, 4, 128'h4030000000000000000000023a4);
sram_add_entry(0, 2, 444, 4, 128'h40300000000000000000000311d);
sram_add_entry(0, 2, 448, 4, 128'h40300000000000000000000995f);
sram_add_entry(0, 2, 452, 4, 128'h403000000000000000000006a35);
sram_add_entry(0, 2, 456, 4, 128'h4030000000000000000000000c8);
sram_add_entry(0, 2, 460, 4, 128'h403000000000000000000003087);
sram_add_entry(0, 2, 464, 4, 128'h40300000000000000000000f1b6);
sram_add_entry(0, 2, 468, 4, 128'h403000000000000000000007805);
sram_add_entry(0, 2, 472, 4, 128'h40300000000000000000000a535);
sram_add_entry(0, 2, 476, 4, 128'h40300000000000000000000ffca);
sram_add_entry(0, 2, 480, 4, 128'h40300000000000000000000fa15);
sram_add_entry(0, 2, 484, 4, 128'h40300000000000000000000de2d);
sram_add_entry(0, 2, 488, 4, 128'h403000000000000000000002fcb);
sram_add_entry(0, 2, 492, 4, 128'h40300000000000000000000432c);
sram_add_entry(0, 2, 496, 4, 128'h40300000000000000000000f151);
sram_add_entry(0, 2, 500, 4, 128'h40300000000000000000000dd1e);
sram_add_entry(0, 2, 504, 4, 128'h40300000000000000000000a8c6);
sram_add_entry(0, 2, 508, 4, 128'h403000000000000000000008146);
sram_add_entry(0, 2, 512, 4, 128'h4030000000000000000000086b9);
sram_add_entry(0, 2, 516, 4, 128'h403000000000000000000006bda);
sram_add_entry(0, 2, 520, 4, 128'h4030000000000000000000035d5);
sram_add_entry(0, 2, 524, 4, 128'h403000000000000000000007354);
sram_add_entry(0, 2, 528, 4, 128'h40300000000000000000000e59b);
sram_add_entry(0, 2, 532, 4, 128'h403000000000000000000004237);
sram_add_entry(0, 2, 536, 4, 128'h403000000000000000000004b8c);
sram_add_entry(0, 2, 540, 4, 128'h403000000000000000000001a7a);
sram_add_entry(0, 2, 544, 4, 128'h40300000000000000000000181b);
sram_add_entry(0, 2, 548, 4, 128'h40300000000000000000000610a);
sram_add_entry(0, 2, 552, 4, 128'h403000000000000000000006087);
sram_add_entry(0, 2, 556, 4, 128'h403000000000000000000005869);
sram_add_entry(0, 2, 560, 4, 128'h403000000000000000000006af7);
sram_add_entry(0, 2, 564, 4, 128'h403000000000000000000009b7f);
sram_add_entry(0, 2, 568, 4, 128'h40300000000000000000000c12a);
sram_add_entry(0, 2, 572, 4, 128'h403000000000000000000007112);
sram_add_entry(0, 2, 576, 4, 128'h40300000000000000000000ff31);
sram_add_entry(0, 2, 580, 4, 128'h40300000000000000000000b651);
sram_add_entry(0, 2, 584, 4, 128'h403000000000000000000004243);
sram_add_entry(0, 2, 588, 4, 128'h40300000000000000000000b299);
sram_add_entry(0, 2, 592, 4, 128'h403000000000000000000007605);
sram_add_entry(0, 2, 596, 4, 128'h40300000000000000000000e4a2);
sram_add_entry(0, 2, 600, 4, 128'h40300000000000000000000e751);
sram_add_entry(0, 2, 604, 4, 128'h40300000000000000000000edf2);
sram_add_entry(0, 2, 608, 4, 128'h403000000000000000000003cfc);
sram_add_entry(0, 2, 612, 4, 128'h40300000000000000000000c7ba);
sram_add_entry(0, 2, 616, 4, 128'h40300000000000000000000c156);
sram_add_entry(0, 2, 620, 4, 128'h4030000000000000000000081aa);
sram_add_entry(0, 2, 624, 4, 128'h40300000000000000000000e58f);
sram_add_entry(0, 2, 628, 4, 128'h403000000000000000000008635);
sram_add_entry(0, 2, 632, 4, 128'h40300000000000000000000af80);
sram_add_entry(0, 2, 636, 4, 128'h40300000000000000000000bad8);
sram_add_entry(0, 2, 640, 4, 128'h40300000000000000000000bcfb);
sram_add_entry(0, 2, 644, 4, 128'h403000000000000000000004b9c);
sram_add_entry(0, 2, 648, 4, 128'h4030000000000000000000072e2);
sram_add_entry(0, 2, 652, 4, 128'h40300000000000000000000c60d);
sram_add_entry(0, 2, 656, 4, 128'h40300000000000000000000a224);
sram_add_entry(0, 2, 660, 4, 128'h40300000000000000000000052f);
sram_add_entry(0, 2, 664, 4, 128'h403000000000000000000001ede);
sram_add_entry(0, 2, 668, 4, 128'h4030000000000000000000041a4);
sram_add_entry(0, 2, 672, 4, 128'h403000000000000000000000615);
sram_add_entry(0, 2, 676, 4, 128'h4030000000000000000000031b1);
sram_add_entry(0, 2, 680, 4, 128'h40300000000000000000000f78f);
sram_add_entry(0, 2, 684, 4, 128'h40300000000000000000000c802);
sram_add_entry(0, 2, 688, 4, 128'h40300000000000000000000829a);
sram_add_entry(0, 2, 692, 4, 128'h403000000000000000000003866);
sram_add_entry(0, 2, 696, 4, 128'h40300000000000000000000e962);
sram_add_entry(0, 2, 700, 4, 128'h40300000000000000000000012f);
sram_add_entry(0, 2, 704, 4, 128'h4030000000000000000000090b9);
sram_add_entry(0, 2, 708, 4, 128'h40300000000000000000000a9bc);
sram_add_entry(0, 2, 712, 4, 128'h403000000000000000000008f6d);
sram_add_entry(0, 2, 716, 4, 128'h40300000000000000000000173a);
sram_add_entry(0, 2, 720, 4, 128'h40300000000000000000000204c);
sram_add_entry(0, 2, 724, 4, 128'h40300000000000000000000f907);
sram_add_entry(0, 2, 728, 4, 128'h40300000000000000000000fc36);
sram_add_entry(0, 2, 732, 4, 128'h40300000000000000000000d4c8);
sram_add_entry(0, 2, 736, 4, 128'h40300000000000000000000cff9);
sram_add_entry(0, 2, 740, 4, 128'h40300000000000000000000167e);
sram_add_entry(0, 2, 744, 4, 128'h40300000000000000000000d549);
sram_add_entry(0, 2, 748, 4, 128'h403000000000000000000000ef1);
sram_add_entry(0, 2, 752, 4, 128'h403000000000000000000000197);
sram_add_entry(0, 2, 756, 4, 128'h40300000000000000000000d74c);
sram_add_entry(0, 2, 760, 4, 128'h40300000000000000000000aa47);
sram_add_entry(0, 2, 764, 4, 128'h40300000000000000000000457b);
sram_add_entry(0, 2, 768, 4, 128'h40300000000000000000000e8d2);
sram_add_entry(0, 2, 772, 4, 128'h4030000000000000000000043db);
sram_add_entry(0, 2, 776, 4, 128'h40300000000000000000000b4cd);
sram_add_entry(0, 2, 780, 4, 128'h403000000000000000000003320);
sram_add_entry(0, 2, 784, 4, 128'h40300000000000000000000f172);
sram_add_entry(0, 2, 788, 4, 128'h40300000000000000000000ab6c);
sram_add_entry(0, 2, 792, 4, 128'h4030000000000000000000010d1);
sram_add_entry(0, 2, 796, 4, 128'h40300000000000000000000c1de);
sram_add_entry(0, 2, 800, 4, 128'h4030000000000000000000004a5);
sram_add_entry(0, 2, 804, 4, 128'h403000000000000000000004677);
sram_add_entry(0, 2, 808, 4, 128'h403000000000000000000001955);
sram_add_entry(0, 2, 812, 4, 128'h403000000000000000000002287);
sram_add_entry(0, 2, 816, 4, 128'h403000000000000000000007fbc);
sram_add_entry(0, 2, 820, 4, 128'h403000000000000000000005226);
sram_add_entry(0, 2, 824, 4, 128'h40300000000000000000000e45e);
sram_add_entry(0, 2, 828, 4, 128'h40300000000000000000000c5d6);
sram_add_entry(0, 2, 832, 4, 128'h40300000000000000000000592e);
sram_add_entry(0, 2, 836, 4, 128'h40300000000000000000000e0dd);
sram_add_entry(0, 2, 840, 4, 128'h403000000000000000000005cd3);
sram_add_entry(0, 2, 844, 4, 128'h403000000000000000000004976);
sram_add_entry(0, 2, 848, 4, 128'h4030000000000000000000055b0);
sram_add_entry(0, 2, 852, 4, 128'h403000000000000000000009ce1);
sram_add_entry(0, 2, 856, 4, 128'h40300000000000000000000981a);
sram_add_entry(0, 2, 860, 4, 128'h40300000000000000000000bc49);
sram_add_entry(0, 2, 864, 4, 128'h403000000000000000000002f11);
sram_add_entry(0, 2, 868, 4, 128'h40300000000000000000000dfe5);
sram_add_entry(0, 2, 872, 4, 128'h40300000000000000000000261b);
sram_add_entry(0, 2, 876, 4, 128'h40300000000000000000000297f);
sram_add_entry(0, 2, 880, 4, 128'h403000000000000000000002d7d);
sram_add_entry(0, 2, 884, 4, 128'h403000000000000000000000ee8);
sram_add_entry(0, 2, 888, 4, 128'h403000000000000000000004561);
sram_add_entry(0, 2, 892, 4, 128'h40300000000000000000000c4c2);
sram_add_entry(0, 2, 896, 4, 128'h40300000000000000000000a32d);
sram_add_entry(0, 2, 900, 4, 128'h40300000000000000000000ff23);
sram_add_entry(0, 2, 904, 4, 128'h40300000000000000000000d60a);
sram_add_entry(0, 2, 908, 4, 128'h403000000000000000000007305);
sram_add_entry(0, 2, 912, 4, 128'h403000000000000000000008bb6);
sram_add_entry(0, 2, 916, 4, 128'h40300000000000000000000ac8c);
sram_add_entry(0, 2, 920, 4, 128'h403000000000000000000008af0);
sram_add_entry(0, 2, 924, 4, 128'h403000000000000000000007c83);
sram_add_entry(0, 2, 928, 4, 128'h40300000000000000000000e1cf);
sram_add_entry(0, 2, 932, 4, 128'h40300000000000000000000e86c);
sram_add_entry(0, 2, 936, 4, 128'h403000000000000000000008c42);
sram_add_entry(0, 2, 940, 4, 128'h4030000000000000000000005f0);
sram_add_entry(0, 2, 944, 4, 128'h403000000000000000000007074);
sram_add_entry(0, 2, 948, 4, 128'h4030000000000000000000014a6);
sram_add_entry(0, 2, 952, 4, 128'h403000000000000000000000576);
sram_add_entry(0, 2, 956, 4, 128'h403000000000000000000005b0b);
sram_add_entry(0, 2, 960, 4, 128'h403000000000000000000004967);
sram_add_entry(0, 2, 964, 4, 128'h4030000000000000000000008e5);
sram_add_entry(0, 2, 968, 4, 128'h403000000000000000000005734);
sram_add_entry(0, 2, 972, 4, 128'h4030000000000000000000077b3);
sram_add_entry(0, 2, 976, 4, 128'h40300000000000000000000de81);
sram_add_entry(0, 2, 980, 4, 128'h403000000000000000000009d79);
sram_add_entry(0, 2, 984, 4, 128'h40300000000000000000000e3fe);
sram_add_entry(0, 2, 988, 4, 128'h403000000000000000000004a66);
sram_add_entry(0, 2, 992, 4, 128'h40300000000000000000000cb9e);
sram_add_entry(0, 2, 996, 4, 128'h403000000000000000000000c1e);
sram_add_entry(0, 2, 1000, 4, 128'h40300000000000000000000da01);
sram_add_entry(0, 2, 1004, 4, 128'h40300000000000000000000fc70);
sram_add_entry(0, 2, 1008, 4, 128'h4030000000000000000000035e4);
sram_add_entry(0, 2, 1012, 4, 128'h403000000000000000000001924);
sram_add_entry(0, 2, 1016, 4, 128'h40300000000000000000000cb60);
sram_add_entry(0, 2, 1020, 4, 128'h403000000000000000000000cb3);
sram_add_entry(0, 2, 1024, 4, 128'h403000000000000000000007107);
sram_add_entry(0, 2, 1028, 4, 128'h40300000000000000000000ef06);
sram_add_entry(0, 2, 1032, 4, 128'h40300000000000000000000b915);
sram_add_entry(0, 2, 1036, 4, 128'h40300000000000000000000569e);
sram_add_entry(0, 2, 1040, 4, 128'h40300000000000000000000a5c6);
sram_add_entry(0, 2, 1044, 4, 128'h403000000000000000000000561);
sram_add_entry(0, 2, 1048, 4, 128'h40300000000000000000000543c);
sram_add_entry(0, 2, 1052, 4, 128'h40300000000000000000000f887);
sram_add_entry(0, 2, 1056, 4, 128'h403000000000000000000002449);
sram_add_entry(0, 2, 1060, 4, 128'h403000000000000000000000aa1);
sram_add_entry(0, 2, 1064, 4, 128'h4030000000000000000000020fc);
sram_add_entry(0, 2, 1068, 4, 128'h4030000000000000000000019c6);
sram_add_entry(0, 2, 1072, 4, 128'h403000000000000000000008d68);
sram_add_entry(0, 2, 1076, 4, 128'h403000000000000000000001fe5);
sram_add_entry(0, 2, 1080, 4, 128'h403000000000000000000008425);
sram_add_entry(0, 2, 1084, 4, 128'h40300000000000000000000ce2c);
sram_add_entry(0, 2, 1088, 4, 128'h403000000000000000000009e07);
sram_add_entry(0, 2, 1092, 4, 128'h40300000000000000000000c360);
sram_add_entry(0, 2, 1096, 4, 128'h4030000000000000000000055a6);
sram_add_entry(0, 2, 1100, 4, 128'h40300000000000000000000d3ce);
sram_add_entry(0, 2, 1104, 4, 128'h4030000000000000000000049ea);
sram_add_entry(0, 2, 1108, 4, 128'h40300000000000000000000e2e3);
sram_add_entry(0, 2, 1112, 4, 128'h403000000000000000000002b4e);
sram_add_entry(0, 2, 1116, 4, 128'h403000000000000000000008ad9);
sram_add_entry(0, 2, 1120, 4, 128'h40300000000000000000000105a);
sram_add_entry(0, 2, 1124, 4, 128'h403000000000000000000000279);
sram_add_entry(0, 2, 1128, 4, 128'h40300000000000000000000933b);
sram_add_entry(0, 2, 1132, 4, 128'h40300000000000000000000a7d8);
sram_add_entry(0, 2, 1136, 4, 128'h403000000000000000000001660);
sram_add_entry(0, 2, 1140, 4, 128'h403000000000000000000002599);
sram_add_entry(0, 2, 1144, 4, 128'h403000000000000000000008360);
sram_add_entry(0, 2, 1148, 4, 128'h403000000000000000000004e54);
sram_add_entry(0, 2, 1152, 4, 128'h403000000000000000000008196);
sram_add_entry(0, 2, 1156, 4, 128'h40300000000000000000000c74f);
sram_add_entry(0, 2, 1160, 4, 128'h40300000000000000000000dbe6);
sram_add_entry(0, 2, 1164, 4, 128'h40300000000000000000000be67);
sram_add_entry(0, 2, 1168, 4, 128'h403000000000000000000003b66);
sram_add_entry(0, 2, 1172, 4, 128'h403000000000000000000000f5d);
sram_add_entry(0, 2, 1176, 4, 128'h403000000000000000000003e97);
sram_add_entry(0, 2, 1180, 4, 128'h4030000000000000000000077cb);
sram_add_entry(0, 2, 1184, 4, 128'h403000000000000000000004ffa);
sram_add_entry(0, 2, 1188, 4, 128'h403000000000000000000005a27);
sram_add_entry(0, 2, 1192, 4, 128'h403000000000000000000004f4a);
sram_add_entry(0, 2, 1196, 4, 128'h40300000000000000000000089b);
sram_add_entry(0, 2, 1200, 4, 128'h40300000000000000000000431f);
sram_add_entry(0, 2, 1204, 4, 128'h40300000000000000000000f164);
sram_add_entry(0, 2, 1208, 4, 128'h40300000000000000000000ae3b);
sram_add_entry(0, 2, 1212, 4, 128'h403000000000000000000004616);
sram_add_entry(0, 2, 1216, 4, 128'h40300000000000000000000e0cf);
sram_add_entry(0, 2, 1220, 4, 128'h403000000000000000000006917);
sram_add_entry(0, 2, 1224, 4, 128'h403000000000000000000002d00);
sram_add_entry(0, 2, 1228, 4, 128'h4030000000000000000000075f9);
sram_add_entry(0, 2, 1232, 4, 128'h403000000000000000000007b29);
sram_add_entry(0, 2, 1236, 4, 128'h4030000000000000000000018be);
sram_add_entry(0, 2, 1240, 4, 128'h4030000000000000000000087d2);
sram_add_entry(0, 2, 1244, 4, 128'h403000000000000000000003974);
sram_add_entry(0, 2, 1248, 4, 128'h4030000000000000000000005c4);
sram_add_entry(0, 2, 1252, 4, 128'h4030000000000000000000018b0);
sram_add_entry(0, 2, 1256, 4, 128'h4030000000000000000000089fd);
sram_add_entry(0, 2, 1260, 4, 128'h403000000000000000000002c4e);
sram_add_entry(0, 2, 1264, 4, 128'h40300000000000000000000417a);
sram_add_entry(0, 2, 1268, 4, 128'h403000000000000000000004888);
sram_add_entry(0, 2, 1272, 4, 128'h403000000000000000000007064);
sram_add_entry(0, 2, 1276, 4, 128'h40300000000000000000000b2bf);
sram_add_entry(0, 2, 1280, 4, 128'h403000000000000000000009d55);
sram_add_entry(0, 2, 1284, 4, 128'h40300000000000000000000ff62);
sram_add_entry(0, 2, 1288, 4, 128'h40300000000000000000000b397);
sram_add_entry(0, 2, 1292, 4, 128'h40300000000000000000000bbdd);
sram_add_entry(0, 2, 1296, 4, 128'h40300000000000000000000871d);
sram_add_entry(0, 2, 1300, 4, 128'h403000000000000000000006fe6);
sram_add_entry(0, 2, 1304, 4, 128'h40300000000000000000000b4f0);
sram_add_entry(0, 2, 1308, 4, 128'h40300000000000000000000343b);
sram_add_entry(0, 2, 1312, 4, 128'h403000000000000000000007848);
sram_add_entry(0, 2, 1316, 4, 128'h40300000000000000000000826c);
sram_add_entry(0, 2, 1320, 4, 128'h40300000000000000000000466e);
sram_add_entry(0, 2, 1324, 4, 128'h403000000000000000000006d50);
sram_add_entry(0, 2, 1328, 4, 128'h40300000000000000000000892d);
sram_add_entry(0, 2, 1332, 4, 128'h403000000000000000000008567);
sram_add_entry(0, 2, 1336, 4, 128'h40300000000000000000000b0d3);
sram_add_entry(0, 2, 1340, 4, 128'h40300000000000000000000c89f);
sram_add_entry(0, 2, 1344, 4, 128'h403000000000000000000002ac3);
sram_add_entry(0, 2, 1348, 4, 128'h403000000000000000000007e5e);
sram_add_entry(0, 2, 1352, 4, 128'h40300000000000000000000d4e5);
sram_add_entry(0, 2, 1356, 4, 128'h40300000000000000000000d1f0);
sram_add_entry(0, 2, 1360, 4, 128'h4030000000000000000000081b0);
sram_add_entry(0, 2, 1364, 4, 128'h40300000000000000000000fcdf);
sram_add_entry(0, 2, 1368, 4, 128'h4030000000000000000000056e8);
sram_add_entry(0, 2, 1372, 4, 128'h403000000000000000000009ba4);
sram_add_entry(0, 2, 1376, 4, 128'h403000000000000000000009667);
sram_add_entry(0, 2, 1380, 4, 128'h403000000000000000000003024);
sram_add_entry(0, 2, 1384, 4, 128'h403000000000000000000000e58);
sram_add_entry(0, 2, 1388, 4, 128'h40300000000000000000000d571);
sram_add_entry(0, 2, 1392, 4, 128'h403000000000000000000007454);
sram_add_entry(0, 2, 1396, 4, 128'h4030000000000000000000011fb);
sram_add_entry(0, 2, 1400, 4, 128'h403000000000000000000006209);
sram_add_entry(0, 2, 1404, 4, 128'h40300000000000000000000e475);
sram_add_entry(0, 2, 1408, 4, 128'h40300000000000000000000c860);
sram_add_entry(0, 2, 1412, 4, 128'h403000000000000000000000781);
sram_add_entry(0, 2, 1416, 4, 128'h403000000000000000000002590);
sram_add_entry(0, 2, 1420, 4, 128'h40300000000000000000000fa8e);
sram_add_entry(0, 2, 1424, 4, 128'h403000000000000000000003f7d);
sram_add_entry(0, 2, 1428, 4, 128'h403000000000000000000000515);
sram_add_entry(0, 2, 1432, 4, 128'h40300000000000000000000b9b3);
sram_add_entry(0, 2, 1436, 4, 128'h403000000000000000000006db1);
sram_add_entry(0, 2, 1440, 4, 128'h40300000000000000000000cde4);
sram_add_entry(0, 2, 1444, 4, 128'h40300000000000000000000ce02);
sram_add_entry(0, 2, 1448, 4, 128'h403000000000000000000004a3c);
sram_add_entry(0, 2, 1452, 4, 128'h403000000000000000000008440);
sram_add_entry(0, 2, 1456, 4, 128'h4030000000000000000000082a7);
sram_add_entry(0, 2, 1460, 4, 128'h40300000000000000000000e481);
sram_add_entry(0, 2, 1464, 4, 128'h403000000000000000000001c1b);
sram_add_entry(0, 2, 1468, 4, 128'h40300000000000000000000819b);
sram_add_entry(0, 2, 1472, 4, 128'h40300000000000000000000e56e);
sram_add_entry(0, 2, 1476, 4, 128'h4030000000000000000000084c7);
sram_add_entry(0, 2, 1480, 4, 128'h403000000000000000000002c16);
sram_add_entry(0, 2, 1484, 4, 128'h403000000000000000000004fb9);
sram_add_entry(0, 2, 1488, 4, 128'h403000000000000000000005dad);
sram_add_entry(0, 2, 1492, 4, 128'h403000000000000000000004e74);
sram_add_entry(0, 2, 1496, 4, 128'h4030000000000000000000030d5);
sram_add_entry(0, 2, 1500, 4, 128'h4030000000000000000000041fa);
sram_add_entry(0, 2, 1504, 4, 128'h40300000000000000000000bf53);
sram_add_entry(0, 2, 1508, 4, 128'h40300000000000000000000901d);
sram_add_entry(0, 2, 1512, 4, 128'h40300000000000000000000f3ee);
sram_add_entry(0, 2, 1516, 4, 128'h403000000000000000000009197);
sram_add_entry(0, 2, 1520, 4, 128'h403000000000000000000001aac);
sram_add_entry(0, 2, 1524, 4, 128'h40300000000000000000000cc69);
sram_add_entry(0, 2, 1528, 4, 128'h403000000000000000000003722);
sram_add_entry(0, 2, 1532, 4, 128'h40300000000000000000000da62);
sram_add_entry(0, 2, 1536, 4, 128'h40300000000000000000000c7f6);
sram_add_entry(0, 2, 1540, 4, 128'h40300000000000000000000e590);
sram_add_entry(0, 2, 1544, 4, 128'h403000000000000000000008354);
sram_add_entry(0, 2, 1548, 4, 128'h40300000000000000000000dee4);
sram_add_entry(0, 2, 1552, 4, 128'h403000000000000000000008a42);
sram_add_entry(0, 2, 1556, 4, 128'h403000000000000000000008249);
sram_add_entry(0, 2, 1560, 4, 128'h40300000000000000000000d7b2);
sram_add_entry(0, 2, 1564, 4, 128'h40300000000000000000000db8d);
sram_add_entry(0, 2, 1568, 4, 128'h403000000000000000000007dca);
sram_add_entry(0, 2, 1572, 4, 128'h403000000000000000000004cb3);
sram_add_entry(0, 2, 1576, 4, 128'h403000000000000000000007648);
sram_add_entry(0, 2, 1580, 4, 128'h4030000000000000000000051a0);
sram_add_entry(0, 2, 1584, 4, 128'h40300000000000000000000fce6);
sram_add_entry(0, 2, 1588, 4, 128'h403000000000000000000001a6e);
sram_add_entry(0, 2, 1592, 4, 128'h403000000000000000000004fab);
sram_add_entry(0, 2, 1596, 4, 128'h40300000000000000000000b664);
sram_add_entry(0, 2, 1600, 4, 128'h403000000000000000000007466);
sram_add_entry(0, 2, 1604, 4, 128'h403000000000000000000005d91);
sram_add_entry(0, 2, 1608, 4, 128'h40300000000000000000000a6d9);
sram_add_entry(0, 2, 1612, 4, 128'h40300000000000000000000066a);
sram_add_entry(0, 2, 1616, 4, 128'h403000000000000000000006c8b);
sram_add_entry(0, 2, 1620, 4, 128'h403000000000000000000007561);
sram_add_entry(0, 2, 1624, 4, 128'h403000000000000000000002b5e);
sram_add_entry(0, 2, 1628, 4, 128'h403000000000000000000005f68);
sram_add_entry(0, 2, 1632, 4, 128'h403000000000000000000008d5a);
sram_add_entry(0, 2, 1636, 4, 128'h403000000000000000000005ff9);
sram_add_entry(0, 2, 1640, 4, 128'h40300000000000000000000aa4a);
sram_add_entry(0, 2, 1644, 4, 128'h403000000000000000000009b48);
sram_add_entry(0, 2, 1648, 4, 128'h40300000000000000000000bab5);
sram_add_entry(0, 2, 1652, 4, 128'h40300000000000000000000e87e);
sram_add_entry(0, 2, 1656, 4, 128'h4030000000000000000000027ff);
sram_add_entry(0, 2, 1660, 4, 128'h40300000000000000000000db49);
sram_add_entry(0, 2, 1664, 4, 128'h40300000000000000000000a716);
sram_add_entry(0, 2, 1668, 4, 128'h40300000000000000000000ea5e);
sram_add_entry(0, 2, 1672, 4, 128'h403000000000000000000009813);
sram_add_entry(0, 2, 1676, 4, 128'h403000000000000000000001c2b);
sram_add_entry(0, 2, 1680, 4, 128'h403000000000000000000005490);
sram_add_entry(0, 2, 1684, 4, 128'h40300000000000000000000dbbc);
sram_add_entry(0, 2, 1688, 4, 128'h40300000000000000000000ba73);
sram_add_entry(0, 2, 1692, 4, 128'h4030000000000000000000022b8);
sram_add_entry(0, 2, 1696, 4, 128'h403000000000000000000004004);
sram_add_entry(0, 2, 1700, 4, 128'h403000000000000000000001d02);
sram_add_entry(0, 2, 1704, 4, 128'h4030000000000000000000032bd);
sram_add_entry(0, 2, 1708, 4, 128'h403000000000000000000005a87);
sram_add_entry(0, 2, 1712, 4, 128'h403000000000000000000001835);
sram_add_entry(0, 2, 1716, 4, 128'h403000000000000000000000348);
sram_add_entry(0, 2, 1720, 4, 128'h403000000000000000000007db8);
sram_add_entry(0, 2, 1724, 4, 128'h4030000000000000000000053a0);
sram_add_entry(0, 2, 1728, 4, 128'h40300000000000000000000094a);
sram_add_entry(0, 2, 1732, 4, 128'h4030000000000000000000068a9);
sram_add_entry(0, 2, 1736, 4, 128'h403000000000000000000006588);
sram_add_entry(0, 2, 1740, 4, 128'h4030000000000000000000054d3);
sram_add_entry(0, 2, 1744, 4, 128'h403000000000000000000007b1e);
sram_add_entry(0, 2, 1748, 4, 128'h403000000000000000000006a07);
sram_add_entry(0, 2, 1752, 4, 128'h40300000000000000000000ecf4);
sram_add_entry(0, 2, 1756, 4, 128'h4030000000000000000000075f1);
sram_add_entry(0, 2, 1760, 4, 128'h4030000000000000000000017b4);
sram_add_entry(0, 2, 1764, 4, 128'h403000000000000000000008fcf);
sram_add_entry(0, 2, 1768, 4, 128'h40300000000000000000000fd38);
sram_add_entry(0, 2, 1772, 4, 128'h4030000000000000000000002d2);
sram_add_entry(0, 2, 1776, 4, 128'h40300000000000000000000c881);
sram_add_entry(0, 2, 1780, 4, 128'h40300000000000000000000bb36);
sram_add_entry(0, 2, 1784, 4, 128'h4030000000000000000000086ff);
sram_add_entry(0, 2, 1788, 4, 128'h40300000000000000000000a23f);
sram_add_entry(0, 2, 1792, 4, 128'h40300000000000000000000d8ec);
sram_add_entry(0, 2, 1796, 4, 128'h403000000000000000000005f93);
sram_add_entry(0, 2, 1800, 4, 128'h403000000000000000000000bc1);
sram_add_entry(0, 2, 1804, 4, 128'h403000000000000000000000144);
sram_add_entry(0, 2, 1808, 4, 128'h40300000000000000000000fdbe);
sram_add_entry(0, 2, 1812, 4, 128'h4030000000000000000000070f4);
sram_add_entry(0, 2, 1816, 4, 128'h403000000000000000000005006);
sram_add_entry(0, 2, 1820, 4, 128'h403000000000000000000004772);
sram_add_entry(0, 2, 1824, 4, 128'h403000000000000000000001aa8);
sram_add_entry(0, 2, 1828, 4, 128'h40300000000000000000000dd72);
sram_add_entry(0, 2, 1832, 4, 128'h403000000000000000000002ec4);
sram_add_entry(0, 2, 1836, 4, 128'h4030000000000000000000033f9);
sram_add_entry(0, 2, 1840, 4, 128'h40300000000000000000000a3f3);
sram_add_entry(0, 2, 1844, 4, 128'h403000000000000000000008144);
sram_add_entry(0, 2, 1848, 4, 128'h403000000000000000000006971);
sram_add_entry(0, 2, 1852, 4, 128'h403000000000000000000003a0f);
sram_add_entry(0, 2, 1856, 4, 128'h40300000000000000000000f3b3);
sram_add_entry(0, 2, 1860, 4, 128'h4030000000000000000000004c3);
sram_add_entry(0, 2, 1864, 4, 128'h4030000000000000000000097a2);
sram_add_entry(0, 2, 1868, 4, 128'h40300000000000000000000191e);
sram_add_entry(0, 2, 1872, 4, 128'h403000000000000000000004c9d);
sram_add_entry(0, 2, 1876, 4, 128'h403000000000000000000001c56);
sram_add_entry(0, 2, 1880, 4, 128'h403000000000000000000004f2e);
sram_add_entry(0, 2, 1884, 4, 128'h403000000000000000000007a32);
sram_add_entry(0, 2, 1888, 4, 128'h40300000000000000000000e58e);
sram_add_entry(0, 2, 1892, 4, 128'h403000000000000000000000fc5);
sram_add_entry(0, 2, 1896, 4, 128'h4030000000000000000000030ab);
sram_add_entry(0, 2, 1900, 4, 128'h403000000000000000000008377);
sram_add_entry(0, 2, 1904, 4, 128'h40300000000000000000000d368);
sram_add_entry(0, 2, 1908, 4, 128'h403000000000000000000006d1d);
sram_add_entry(0, 2, 1912, 4, 128'h4030000000000000000000023a3);
sram_add_entry(0, 2, 1916, 4, 128'h403000000000000000000004845);
sram_add_entry(0, 2, 1920, 4, 128'h40300000000000000000000992e);
sram_add_entry(0, 2, 1924, 4, 128'h403000000000000000000009aad);
sram_add_entry(0, 2, 1928, 4, 128'h403000000000000000000000c17);
sram_add_entry(0, 2, 1932, 4, 128'h40300000000000000000000ce74);
sram_add_entry(0, 2, 1936, 4, 128'h40300000000000000000000a3bc);
sram_add_entry(0, 2, 1940, 4, 128'h40300000000000000000000af3e);
sram_add_entry(0, 2, 1944, 4, 128'h40300000000000000000000f44a);
sram_add_entry(0, 2, 1948, 4, 128'h40300000000000000000000abdc);
sram_add_entry(0, 2, 1952, 4, 128'h403000000000000000000001ffa);
sram_add_entry(0, 2, 1956, 4, 128'h40300000000000000000000bbe8);
sram_add_entry(0, 2, 1960, 4, 128'h40300000000000000000000ce02);
sram_add_entry(0, 2, 1964, 4, 128'h403000000000000000000000f7a);
sram_add_entry(0, 2, 1968, 4, 128'h403000000000000000000000b92);
sram_add_entry(0, 2, 1972, 4, 128'h40300000000000000000000371a);
sram_add_entry(0, 2, 1976, 4, 128'h403000000000000000000005154);
sram_add_entry(0, 2, 1980, 4, 128'h40300000000000000000000244d);
sram_add_entry(0, 2, 1984, 4, 128'h40300000000000000000000d841);
sram_add_entry(0, 2, 1988, 4, 128'h403000000000000000000007799);
sram_add_entry(0, 2, 1992, 4, 128'h403000000000000000000004853);
sram_add_entry(0, 2, 1996, 4, 128'h403000000000000000000009615);
sram_add_entry(0, 2, 2000, 4, 128'h4030000000000000000000025af);
sram_add_entry(0, 2, 2004, 4, 128'h4030000000000000000000025f9);
sram_add_entry(0, 2, 2008, 4, 128'h403000000000000000000002c36);
sram_add_entry(0, 2, 2012, 4, 128'h403000000000000000000006575);
sram_add_entry(0, 2, 2016, 4, 128'h403000000000000000000003684);
sram_add_entry(0, 2, 2020, 4, 128'h40300000000000000000000f639);
sram_add_entry(0, 2, 2024, 4, 128'h4030000000000000000000026d1);
sram_add_entry(0, 2, 2028, 4, 128'h4030000000000000000000013dd);
sram_add_entry(0, 2, 2032, 4, 128'h403000000000000000000003335);
sram_add_entry(0, 2, 2036, 4, 128'h40300000000000000000000e6ea);
sram_add_entry(0, 2, 2040, 4, 128'h403000000000000000000001403);
sram_add_entry(0, 2, 2044, 4, 128'h40300000000000000000000b48a);
sram_add_entry(0, 2, 2048, 4, 128'h403000000000000000000003a1b);
sram_add_entry(0, 2, 2052, 4, 128'h40300000000000000000000c0f4);
sram_add_entry(0, 2, 2056, 4, 128'h40300000000000000000000b6f5);
sram_add_entry(0, 2, 2060, 4, 128'h403000000000000000000005c2f);
sram_add_entry(0, 2, 2064, 4, 128'h4030000000000000000000062e1);
sram_add_entry(0, 2, 2068, 4, 128'h40300000000000000000000c121);
sram_add_entry(0, 2, 2072, 4, 128'h40300000000000000000000c629);
sram_add_entry(0, 2, 2076, 4, 128'h4030000000000000000000019d2);
sram_add_entry(0, 2, 2080, 4, 128'h403000000000000000000009600);
sram_add_entry(0, 2, 2084, 4, 128'h403000000000000000000000b54);
sram_add_entry(0, 2, 2088, 4, 128'h40300000000000000000000d9db);
sram_add_entry(0, 2, 2092, 4, 128'h40300000000000000000000284a);
sram_add_entry(0, 2, 2096, 4, 128'h403000000000000000000006511);
sram_add_entry(0, 2, 2100, 4, 128'h40300000000000000000000b42e);
sram_add_entry(0, 2, 2104, 4, 128'h40300000000000000000000a05a);
sram_add_entry(0, 2, 2108, 4, 128'h403000000000000000000004f13);
sram_add_entry(0, 2, 2112, 4, 128'h4030000000000000000000005ae);
sram_add_entry(0, 2, 2116, 4, 128'h403000000000000000000002d8c);
sram_add_entry(0, 2, 2120, 4, 128'h403000000000000000000002bff);
sram_add_entry(0, 2, 2124, 4, 128'h403000000000000000000009abe);
sram_add_entry(0, 2, 2128, 4, 128'h40300000000000000000000cfd9);
sram_add_entry(0, 2, 2132, 4, 128'h403000000000000000000003957);
sram_add_entry(0, 2, 2136, 4, 128'h403000000000000000000004efb);
sram_add_entry(0, 2, 2140, 4, 128'h40300000000000000000000dd5e);
sram_add_entry(0, 2, 2144, 4, 128'h40300000000000000000000800e);
sram_add_entry(0, 2, 2148, 4, 128'h403000000000000000000001697);
sram_add_entry(0, 2, 2152, 4, 128'h4030000000000000000000042ce);
sram_add_entry(0, 2, 2156, 4, 128'h40300000000000000000000bcbf);
sram_add_entry(0, 2, 2160, 4, 128'h403000000000000000000008541);
sram_add_entry(0, 2, 2164, 4, 128'h4030000000000000000000085d1);
sram_add_entry(0, 2, 2168, 4, 128'h403000000000000000000003385);
sram_add_entry(0, 2, 2172, 4, 128'h40300000000000000000000708c);
sram_add_entry(0, 2, 2176, 4, 128'h403000000000000000000002082);
sram_add_entry(0, 2, 2180, 4, 128'h40300000000000000000000055b);
sram_add_entry(0, 2, 2184, 4, 128'h4030000000000000000000015db);
sram_add_entry(0, 2, 2188, 4, 128'h40300000000000000000000614f);
sram_add_entry(0, 2, 2192, 4, 128'h4030000000000000000000013b4);
sram_add_entry(0, 2, 2196, 4, 128'h403000000000000000000004a8b);
sram_add_entry(0, 2, 2200, 4, 128'h40300000000000000000000d328);
sram_add_entry(0, 2, 2204, 4, 128'h403000000000000000000002219);
sram_add_entry(0, 2, 2208, 4, 128'h40300000000000000000000fdef);
sram_add_entry(0, 2, 2212, 4, 128'h40300000000000000000000cab1);
sram_add_entry(0, 2, 2216, 4, 128'h403000000000000000000008dc9);
sram_add_entry(0, 2, 2220, 4, 128'h403000000000000000000008a3e);
sram_add_entry(0, 2, 2224, 4, 128'h403000000000000000000002949);
sram_add_entry(0, 2, 2228, 4, 128'h40300000000000000000000d515);
sram_add_entry(0, 2, 2232, 4, 128'h40300000000000000000000a7ab);
sram_add_entry(0, 2, 2236, 4, 128'h403000000000000000000008155);
sram_add_entry(0, 2, 2240, 4, 128'h40300000000000000000000bbc5);
sram_add_entry(0, 2, 2244, 4, 128'h403000000000000000000005035);
sram_add_entry(0, 2, 2248, 4, 128'h40300000000000000000000b93f);
sram_add_entry(0, 2, 2252, 4, 128'h4030000000000000000000037bb);
sram_add_entry(0, 2, 2256, 4, 128'h403000000000000000000006387);
sram_add_entry(0, 2, 2260, 4, 128'h40300000000000000000000338f);
sram_add_entry(0, 2, 2264, 4, 128'h4030000000000000000000026a6);
sram_add_entry(0, 2, 2268, 4, 128'h40300000000000000000000206d);
sram_add_entry(0, 2, 2272, 4, 128'h403000000000000000000008535);
sram_add_entry(0, 2, 2276, 4, 128'h403000000000000000000001b88);
sram_add_entry(0, 2, 2280, 4, 128'h40300000000000000000000fbe6);
sram_add_entry(0, 2, 2284, 4, 128'h40300000000000000000000e4bf);
sram_add_entry(0, 2, 2288, 4, 128'h40300000000000000000000a5a6);
sram_add_entry(0, 2, 2292, 4, 128'h403000000000000000000009f00);
sram_add_entry(0, 2, 2296, 4, 128'h403000000000000000000006530);
sram_add_entry(0, 2, 2300, 4, 128'h4030000000000000000000037d5);
sram_add_entry(0, 2, 2304, 4, 128'h403000000000000000000009b09);
sram_add_entry(0, 2, 2308, 4, 128'h40300000000000000000000a8bd);
sram_add_entry(0, 2, 2312, 4, 128'h40300000000000000000000e4f1);
sram_add_entry(0, 2, 2316, 4, 128'h40300000000000000000000d34e);
sram_add_entry(0, 2, 2320, 4, 128'h4030000000000000000000028f9);
sram_add_entry(0, 2, 2324, 4, 128'h403000000000000000000007c60);
sram_add_entry(0, 2, 2328, 4, 128'h40300000000000000000000d4d5);
sram_add_entry(0, 2, 2332, 4, 128'h403000000000000000000004278);
sram_add_entry(0, 2, 2336, 4, 128'h403000000000000000000002823);
sram_add_entry(0, 2, 2340, 4, 128'h40300000000000000000000df68);
sram_add_entry(0, 2, 2344, 4, 128'h403000000000000000000007947);
sram_add_entry(0, 2, 2348, 4, 128'h40300000000000000000000a587);
sram_add_entry(0, 2, 2352, 4, 128'h4030000000000000000000051ce);
sram_add_entry(0, 2, 2356, 4, 128'h40300000000000000000000110a);
sram_add_entry(0, 2, 2360, 4, 128'h40300000000000000000000effe);
sram_add_entry(0, 2, 2364, 4, 128'h403000000000000000000000d97);
sram_add_entry(0, 2, 2368, 4, 128'h403000000000000000000002191);
sram_add_entry(0, 2, 2372, 4, 128'h40300000000000000000000a878);
sram_add_entry(0, 2, 2376, 4, 128'h40300000000000000000000f873);
sram_add_entry(0, 2, 2380, 4, 128'h40300000000000000000000df00);
sram_add_entry(0, 2, 2384, 4, 128'h403000000000000000000008139);
sram_add_entry(0, 2, 2388, 4, 128'h403000000000000000000005538);
sram_add_entry(0, 2, 2392, 4, 128'h40300000000000000000000e1ce);
sram_add_entry(0, 2, 2396, 4, 128'h4030000000000000000000034dc);
sram_add_entry(0, 2, 2400, 4, 128'h40300000000000000000000751e);
sram_add_entry(0, 2, 2404, 4, 128'h4030000000000000000000048e3);
sram_add_entry(0, 2, 2408, 4, 128'h40300000000000000000000d719);
sram_add_entry(0, 2, 2412, 4, 128'h403000000000000000000006f67);
sram_add_entry(0, 2, 2416, 4, 128'h40300000000000000000000d5af);
sram_add_entry(0, 2, 2420, 4, 128'h403000000000000000000001c7c);
sram_add_entry(0, 2, 2424, 4, 128'h403000000000000000000005a36);
sram_add_entry(0, 2, 2428, 4, 128'h403000000000000000000005647);
sram_add_entry(0, 2, 2432, 4, 128'h40300000000000000000000a79e);
sram_add_entry(0, 2, 2436, 4, 128'h40300000000000000000000b278);
sram_add_entry(0, 2, 2440, 4, 128'h4030000000000000000000040bf);
sram_add_entry(0, 2, 2444, 4, 128'h40300000000000000000000799e);
sram_add_entry(0, 2, 2448, 4, 128'h40300000000000000000000b51c);
sram_add_entry(0, 2, 2452, 4, 128'h40300000000000000000000eb9a);
sram_add_entry(0, 2, 2456, 4, 128'h403000000000000000000003e44);
sram_add_entry(0, 2, 2460, 4, 128'h4030000000000000000000088bd);
sram_add_entry(0, 2, 2464, 4, 128'h403000000000000000000006126);
sram_add_entry(0, 2, 2468, 4, 128'h40300000000000000000000e67b);
sram_add_entry(0, 2, 2472, 4, 128'h40300000000000000000000b998);
sram_add_entry(0, 2, 2476, 4, 128'h4030000000000000000000082fe);
sram_add_entry(0, 2, 2480, 4, 128'h403000000000000000000003203);
sram_add_entry(0, 2, 2484, 4, 128'h40300000000000000000000d92b);
sram_add_entry(0, 2, 2488, 4, 128'h4030000000000000000000080ec);
sram_add_entry(0, 2, 2492, 4, 128'h403000000000000000000007aa1);
sram_add_entry(0, 2, 2496, 4, 128'h40300000000000000000000fff3);
sram_add_entry(0, 2, 2500, 4, 128'h4030000000000000000000019f1);
sram_add_entry(0, 2, 2504, 4, 128'h40300000000000000000000e2d3);
sram_add_entry(0, 2, 2508, 4, 128'h403000000000000000000001c4b);
sram_add_entry(0, 2, 2512, 4, 128'h40300000000000000000000f785);
sram_add_entry(0, 2, 2516, 4, 128'h403000000000000000000006e92);
sram_add_entry(0, 2, 2520, 4, 128'h403000000000000000000008164);
sram_add_entry(0, 2, 2524, 4, 128'h40300000000000000000000c136);
sram_add_entry(0, 2, 2528, 4, 128'h4030000000000000000000079d2);
sram_add_entry(0, 2, 2532, 4, 128'h40300000000000000000000e175);
sram_add_entry(0, 2, 2536, 4, 128'h403000000000000000000006eda);
sram_add_entry(0, 2, 2540, 4, 128'h403000000000000000000006c68);
sram_add_entry(0, 2, 2544, 4, 128'h40300000000000000000000be89);
sram_add_entry(0, 2, 2548, 4, 128'h40300000000000000000000d49f);
sram_add_entry(0, 2, 2552, 4, 128'h403000000000000000000009a7f);
sram_add_entry(0, 2, 2556, 4, 128'h403000000000000000000004960);
sram_add_entry(0, 2, 2560, 4, 128'h403000000000000000000001bc1);
sram_add_entry(0, 2, 2564, 4, 128'h40300000000000000000000144e);
sram_add_entry(0, 2, 2568, 4, 128'h40300000000000000000000779c);
sram_add_entry(0, 2, 2572, 4, 128'h40300000000000000000000871a);
sram_add_entry(0, 2, 2576, 4, 128'h403000000000000000000001b85);
sram_add_entry(0, 2, 2580, 4, 128'h403000000000000000000000b1e);
sram_add_entry(0, 2, 2584, 4, 128'h40300000000000000000000573c);
sram_add_entry(0, 2, 2588, 4, 128'h4030000000000000000000043ec);
sram_add_entry(0, 2, 2592, 4, 128'h403000000000000000000009e70);
sram_add_entry(0, 2, 2596, 4, 128'h403000000000000000000007bbb);
sram_add_entry(0, 2, 2600, 4, 128'h4030000000000000000000058a8);
sram_add_entry(0, 2, 2604, 4, 128'h40300000000000000000000bb95);
sram_add_entry(0, 2, 2608, 4, 128'h403000000000000000000004ee1);
sram_add_entry(0, 2, 2612, 4, 128'h40300000000000000000000cd5e);
sram_add_entry(0, 2, 2616, 4, 128'h40300000000000000000000855f);
sram_add_entry(0, 2, 2620, 4, 128'h403000000000000000000007a49);
sram_add_entry(0, 2, 2624, 4, 128'h403000000000000000000001c06);
sram_add_entry(0, 2, 2628, 4, 128'h40300000000000000000000dc16);
sram_add_entry(0, 2, 2632, 4, 128'h40300000000000000000000618d);
sram_add_entry(0, 2, 2636, 4, 128'h403000000000000000000007ea0);
sram_add_entry(0, 2, 2640, 4, 128'h40300000000000000000000d910);
sram_add_entry(0, 2, 2644, 4, 128'h40300000000000000000000dc31);
sram_add_entry(0, 2, 2648, 4, 128'h4030000000000000000000088aa);
sram_add_entry(0, 2, 2652, 4, 128'h4030000000000000000000089fe);
sram_add_entry(0, 2, 2656, 4, 128'h40300000000000000000000f777);
sram_add_entry(0, 2, 2660, 4, 128'h4030000000000000000000028d5);
sram_add_entry(0, 2, 2664, 4, 128'h403000000000000000000005497);
sram_add_entry(0, 2, 2668, 4, 128'h403000000000000000000009db1);
sram_add_entry(0, 2, 2672, 4, 128'h403000000000000000000000570);
sram_add_entry(0, 2, 2676, 4, 128'h40300000000000000000000e79a);
sram_add_entry(0, 2, 2680, 4, 128'h40300000000000000000000aa71);
sram_add_entry(0, 2, 2684, 4, 128'h40300000000000000000000dd36);
sram_add_entry(0, 2, 2688, 4, 128'h4030000000000000000000077a3);
sram_add_entry(0, 2, 2692, 4, 128'h403000000000000000000002946);
sram_add_entry(0, 2, 2696, 4, 128'h40300000000000000000000c3d1);
sram_add_entry(0, 2, 2700, 4, 128'h40300000000000000000000884e);
sram_add_entry(0, 2, 2704, 4, 128'h40300000000000000000000552c);
sram_add_entry(0, 2, 2708, 4, 128'h40300000000000000000000418f);
sram_add_entry(0, 2, 2712, 4, 128'h4030000000000000000000002d0);
sram_add_entry(0, 2, 2716, 4, 128'h403000000000000000000001688);
sram_add_entry(0, 2, 2720, 4, 128'h40300000000000000000000d1ea);
sram_add_entry(0, 2, 2724, 4, 128'h40300000000000000000000ed72);
sram_add_entry(0, 2, 2728, 4, 128'h403000000000000000000004b54);
sram_add_entry(0, 2, 2732, 4, 128'h40300000000000000000000a5ad);
sram_add_entry(0, 2, 2736, 4, 128'h403000000000000000000002270);
sram_add_entry(0, 2, 2740, 4, 128'h403000000000000000000007c75);
sram_add_entry(0, 2, 2744, 4, 128'h403000000000000000000003d8c);
sram_add_entry(0, 2, 2748, 4, 128'h4030000000000000000000054cc);
sram_add_entry(0, 2, 2752, 4, 128'h403000000000000000000008f89);
sram_add_entry(0, 2, 2756, 4, 128'h40300000000000000000000641e);
sram_add_entry(0, 2, 2760, 4, 128'h40300000000000000000000066d);
sram_add_entry(0, 2, 2764, 4, 128'h40300000000000000000000f56a);
sram_add_entry(0, 2, 2768, 4, 128'h403000000000000000000000478);
sram_add_entry(0, 2, 2772, 4, 128'h40300000000000000000000668d);
sram_add_entry(0, 2, 2776, 4, 128'h40300000000000000000000a161);
sram_add_entry(0, 2, 2780, 4, 128'h403000000000000000000006b35);
sram_add_entry(0, 2, 2784, 4, 128'h403000000000000000000005b97);
sram_add_entry(0, 2, 2788, 4, 128'h40300000000000000000000f63c);
sram_add_entry(0, 2, 2792, 4, 128'h403000000000000000000005629);
sram_add_entry(0, 2, 2796, 4, 128'h403000000000000000000002745);
sram_add_entry(0, 2, 2800, 4, 128'h40300000000000000000000232e);
sram_add_entry(0, 4, 0, 4, 128'h7ab000000000000000000deadbf);
sram_add_entry(0, 4, 4, 4, 128'h403000000000000000000006814);
sram_add_entry(0, 4, 8, 4, 128'h40300000000000000000000c070);
sram_add_entry(0, 4, 12, 4, 128'h403000000000000000000009740);
sram_add_entry(0, 4, 16, 4, 128'h40300000000000000000000c6fc);
sram_add_entry(0, 4, 20, 4, 128'h40300000000000000000000123a);
sram_add_entry(0, 4, 24, 4, 128'h403000000000000000000007780);
sram_add_entry(0, 4, 28, 4, 128'h40300000000000000000000a3a1);
sram_add_entry(0, 4, 32, 4, 128'h403000000000000000000003259);
sram_add_entry(0, 4, 36, 4, 128'h40300000000000000000000b3e9);
sram_add_entry(0, 4, 40, 4, 128'h403000000000000000000006bec);
sram_add_entry(0, 4, 44, 4, 128'h403000000000000000000003843);
sram_add_entry(0, 4, 48, 4, 128'h4030000000000000000000089af);
sram_add_entry(0, 4, 52, 4, 128'h403000000000000000000008c78);
sram_add_entry(0, 4, 56, 4, 128'h4030000000000000000000018e7);
sram_add_entry(0, 4, 60, 4, 128'h4030000000000000000000075ae);
sram_add_entry(0, 4, 64, 4, 128'h4030000000000000000000080c5);
sram_add_entry(0, 4, 68, 4, 128'h403000000000000000000009a32);
sram_add_entry(0, 4, 72, 4, 128'h40300000000000000000000e7a9);
sram_add_entry(0, 4, 76, 4, 128'h40300000000000000000000ebf7);
sram_add_entry(0, 4, 80, 4, 128'h40300000000000000000000cd9a);
sram_add_entry(0, 4, 84, 4, 128'h403000000000000000000002365);
sram_add_entry(0, 4, 88, 4, 128'h403000000000000000000009688);
sram_add_entry(0, 4, 92, 4, 128'h40300000000000000000000e859);
sram_add_entry(0, 4, 96, 4, 128'h40300000000000000000000b77b);
sram_add_entry(0, 4, 100, 4, 128'h403000000000000000000002430);
sram_add_entry(0, 4, 104, 4, 128'h40300000000000000000000cb20);
sram_add_entry(0, 4, 108, 4, 128'h40300000000000000000000a1e3);
sram_add_entry(0, 4, 112, 4, 128'h403000000000000000000000acc);
sram_add_entry(0, 4, 116, 4, 128'h40300000000000000000000eb72);
sram_add_entry(0, 4, 120, 4, 128'h403000000000000000000000f78);
sram_add_entry(0, 4, 124, 4, 128'h403000000000000000000007d85);
sram_add_entry(0, 4, 128, 4, 128'h40300000000000000000000d586);
sram_add_entry(0, 4, 132, 4, 128'h403000000000000000000007dab);
sram_add_entry(0, 4, 136, 4, 128'h40300000000000000000000cb04);
sram_add_entry(0, 4, 140, 4, 128'h403000000000000000000009cbc);
sram_add_entry(0, 4, 144, 4, 128'h40300000000000000000000e211);
sram_add_entry(0, 4, 148, 4, 128'h40300000000000000000000b146);
sram_add_entry(0, 4, 152, 4, 128'h403000000000000000000004e87);
sram_add_entry(0, 4, 156, 4, 128'h40300000000000000000000597c);
sram_add_entry(0, 4, 160, 4, 128'h403000000000000000000003e12);
sram_add_entry(0, 4, 164, 4, 128'h403000000000000000000009949);
sram_add_entry(0, 4, 168, 4, 128'h4030000000000000000000094fa);
sram_add_entry(0, 4, 172, 4, 128'h40300000000000000000000cdb2);
sram_add_entry(0, 4, 176, 4, 128'h40300000000000000000000fe66);
sram_add_entry(0, 4, 180, 4, 128'h40300000000000000000000c0c2);
sram_add_entry(0, 4, 184, 4, 128'h40300000000000000000000f232);
sram_add_entry(0, 4, 188, 4, 128'h40300000000000000000000a7be);
sram_add_entry(0, 4, 192, 4, 128'h403000000000000000000000fcd);
sram_add_entry(0, 4, 196, 4, 128'h40300000000000000000000b422);
sram_add_entry(0, 4, 200, 4, 128'h40300000000000000000000d35e);
sram_add_entry(0, 4, 204, 4, 128'h40300000000000000000000a927);
sram_add_entry(0, 4, 208, 4, 128'h40300000000000000000000b0b8);
sram_add_entry(0, 4, 212, 4, 128'h403000000000000000000006f6b);
sram_add_entry(0, 4, 216, 4, 128'h40300000000000000000000bd1d);
sram_add_entry(0, 4, 220, 4, 128'h40300000000000000000000981d);
sram_add_entry(0, 4, 224, 4, 128'h403000000000000000000000afd);
sram_add_entry(0, 4, 228, 4, 128'h40300000000000000000000dd25);
sram_add_entry(0, 4, 232, 4, 128'h403000000000000000000006dac);
sram_add_entry(0, 4, 236, 4, 128'h4030000000000000000000025d5);
sram_add_entry(0, 4, 240, 4, 128'h403000000000000000000005737);
sram_add_entry(0, 4, 244, 4, 128'h40300000000000000000000964f);
sram_add_entry(0, 4, 248, 4, 128'h40300000000000000000000ee96);
sram_add_entry(0, 4, 252, 4, 128'h403000000000000000000008464);
sram_add_entry(0, 4, 256, 4, 128'h40300000000000000000000be76);
sram_add_entry(0, 4, 260, 4, 128'h403000000000000000000005a21);
sram_add_entry(0, 4, 264, 4, 128'h40300000000000000000000550d);
sram_add_entry(0, 4, 268, 4, 128'h40300000000000000000000ebb4);
sram_add_entry(0, 4, 272, 4, 128'h40300000000000000000000cc55);
sram_add_entry(0, 4, 276, 4, 128'h403000000000000000000007a15);
sram_add_entry(0, 4, 280, 4, 128'h40300000000000000000000d887);
sram_add_entry(0, 4, 284, 4, 128'h403000000000000000000006379);
sram_add_entry(0, 4, 288, 4, 128'h40300000000000000000000843c);
sram_add_entry(0, 4, 292, 4, 128'h40300000000000000000000353c);
sram_add_entry(0, 4, 296, 4, 128'h4030000000000000000000043e1);
sram_add_entry(0, 4, 300, 4, 128'h403000000000000000000009c19);
sram_add_entry(0, 4, 304, 4, 128'h40300000000000000000000cd0b);
sram_add_entry(0, 4, 308, 4, 128'h403000000000000000000005254);
sram_add_entry(0, 4, 312, 4, 128'h40300000000000000000000d8e8);
sram_add_entry(0, 4, 316, 4, 128'h40300000000000000000000e7a6);
sram_add_entry(0, 4, 320, 4, 128'h40300000000000000000000a32f);
sram_add_entry(0, 4, 324, 4, 128'h40300000000000000000000fb8d);
sram_add_entry(0, 4, 328, 4, 128'h4030000000000000000000039f9);
sram_add_entry(0, 4, 332, 4, 128'h403000000000000000000007d79);
sram_add_entry(0, 4, 336, 4, 128'h40300000000000000000000b263);
sram_add_entry(0, 4, 340, 4, 128'h40300000000000000000000b28d);
sram_add_entry(0, 4, 344, 4, 128'h403000000000000000000005639);
sram_add_entry(0, 4, 348, 4, 128'h403000000000000000000002011);
sram_add_entry(0, 4, 352, 4, 128'h40300000000000000000000bf31);
sram_add_entry(0, 4, 356, 4, 128'h40300000000000000000000902b);
sram_add_entry(0, 4, 360, 4, 128'h40300000000000000000000889d);
sram_add_entry(0, 4, 364, 4, 128'h403000000000000000000001e7e);
sram_add_entry(0, 4, 368, 4, 128'h4030000000000000000000066b7);
sram_add_entry(0, 4, 372, 4, 128'h40300000000000000000000e7a4);
sram_add_entry(0, 4, 376, 4, 128'h40300000000000000000000f191);
sram_add_entry(0, 4, 380, 4, 128'h40300000000000000000000a000);
sram_add_entry(0, 4, 384, 4, 128'h40300000000000000000000304f);
sram_add_entry(0, 4, 388, 4, 128'h40300000000000000000000cc62);
sram_add_entry(0, 4, 392, 4, 128'h4030000000000000000000042cd);
sram_add_entry(0, 4, 396, 4, 128'h40300000000000000000000b26a);
sram_add_entry(0, 4, 400, 4, 128'h40300000000000000000000c7be);
sram_add_entry(0, 4, 404, 4, 128'h40300000000000000000000b1b8);
sram_add_entry(0, 4, 408, 4, 128'h40300000000000000000000fac7);
sram_add_entry(0, 4, 412, 4, 128'h4030000000000000000000022e7);
sram_add_entry(0, 4, 416, 4, 128'h40300000000000000000000085e);
sram_add_entry(0, 4, 420, 4, 128'h403000000000000000000006156);
sram_add_entry(0, 4, 424, 4, 128'h403000000000000000000004e18);
sram_add_entry(0, 4, 428, 4, 128'h403000000000000000000008df4);
sram_add_entry(0, 4, 432, 4, 128'h40300000000000000000000c184);
sram_add_entry(0, 4, 436, 4, 128'h4030000000000000000000024f9);
sram_add_entry(0, 4, 440, 4, 128'h4030000000000000000000055a9);
sram_add_entry(0, 4, 444, 4, 128'h403000000000000000000007d2c);
sram_add_entry(0, 4, 448, 4, 128'h403000000000000000000008b7b);
sram_add_entry(0, 4, 452, 4, 128'h403000000000000000000006e62);
sram_add_entry(0, 4, 456, 4, 128'h40300000000000000000000aa01);
sram_add_entry(0, 4, 460, 4, 128'h40300000000000000000000b523);
sram_add_entry(0, 4, 464, 4, 128'h403000000000000000000009dba);
sram_add_entry(0, 4, 468, 4, 128'h40300000000000000000000c4e7);
sram_add_entry(0, 4, 472, 4, 128'h40300000000000000000000df70);
sram_add_entry(0, 4, 476, 4, 128'h403000000000000000000000a6b);
sram_add_entry(0, 4, 480, 4, 128'h403000000000000000000003efb);
sram_add_entry(0, 4, 484, 4, 128'h40300000000000000000000c13b);
sram_add_entry(0, 4, 488, 4, 128'h40300000000000000000000dd53);
sram_add_entry(0, 4, 492, 4, 128'h40300000000000000000000dc42);
sram_add_entry(0, 4, 496, 4, 128'h40300000000000000000000d019);
sram_add_entry(0, 4, 500, 4, 128'h403000000000000000000004ac7);
sram_add_entry(0, 4, 504, 4, 128'h403000000000000000000001c65);
sram_add_entry(0, 4, 508, 4, 128'h40300000000000000000000c12e);
sram_add_entry(0, 4, 512, 4, 128'h403000000000000000000006cc2);
sram_add_entry(0, 4, 516, 4, 128'h403000000000000000000001979);
sram_add_entry(0, 4, 520, 4, 128'h403000000000000000000003003);
sram_add_entry(0, 4, 524, 4, 128'h40300000000000000000000e7fc);
sram_add_entry(0, 4, 528, 4, 128'h40300000000000000000000b67b);
sram_add_entry(0, 4, 532, 4, 128'h40300000000000000000000d14d);
sram_add_entry(0, 4, 536, 4, 128'h403000000000000000000008684);
sram_add_entry(0, 4, 540, 4, 128'h403000000000000000000006940);
sram_add_entry(0, 4, 544, 4, 128'h4030000000000000000000034fd);
sram_add_entry(0, 4, 548, 4, 128'h4030000000000000000000089e2);
sram_add_entry(0, 4, 552, 4, 128'h40300000000000000000000da12);
sram_add_entry(0, 4, 556, 4, 128'h403000000000000000000000864);
sram_add_entry(0, 4, 560, 4, 128'h40300000000000000000000b1ee);
sram_add_entry(0, 4, 564, 4, 128'h40300000000000000000000b1e4);
sram_add_entry(0, 4, 568, 4, 128'h40300000000000000000000cc72);
sram_add_entry(0, 4, 572, 4, 128'h40300000000000000000000be14);
sram_add_entry(0, 4, 576, 4, 128'h40300000000000000000000cda4);
sram_add_entry(0, 4, 580, 4, 128'h4030000000000000000000040c1);
sram_add_entry(0, 4, 584, 4, 128'h403000000000000000000005d6d);
sram_add_entry(0, 4, 588, 4, 128'h403000000000000000000004fc3);
sram_add_entry(0, 4, 592, 4, 128'h40300000000000000000000c62b);
sram_add_entry(0, 4, 596, 4, 128'h40300000000000000000000f641);
sram_add_entry(0, 4, 600, 4, 128'h40300000000000000000000cef3);
sram_add_entry(0, 4, 604, 4, 128'h403000000000000000000000585);
sram_add_entry(0, 4, 608, 4, 128'h40300000000000000000000058e);
sram_add_entry(0, 4, 612, 4, 128'h403000000000000000000008895);
sram_add_entry(0, 4, 616, 4, 128'h403000000000000000000008e73);
sram_add_entry(0, 4, 620, 4, 128'h40300000000000000000000bc7d);
sram_add_entry(0, 4, 624, 4, 128'h403000000000000000000000d48);
sram_add_entry(0, 4, 628, 4, 128'h40300000000000000000000de40);
sram_add_entry(0, 4, 632, 4, 128'h403000000000000000000000c40);
sram_add_entry(0, 4, 636, 4, 128'h40300000000000000000000200d);
sram_add_entry(0, 4, 640, 4, 128'h403000000000000000000001ac3);
sram_add_entry(0, 4, 644, 4, 128'h403000000000000000000007006);
sram_add_entry(0, 4, 648, 4, 128'h40300000000000000000000bc2d);
sram_add_entry(0, 4, 652, 4, 128'h40300000000000000000000da27);
sram_add_entry(0, 4, 656, 4, 128'h40300000000000000000000e8d9);
sram_add_entry(0, 4, 660, 4, 128'h40300000000000000000000cf50);
sram_add_entry(0, 4, 664, 4, 128'h4030000000000000000000053d6);
sram_add_entry(0, 4, 668, 4, 128'h403000000000000000000008515);
sram_add_entry(0, 4, 672, 4, 128'h403000000000000000000003f78);
sram_add_entry(0, 4, 676, 4, 128'h40300000000000000000000f457);
sram_add_entry(0, 4, 680, 4, 128'h4030000000000000000000044bc);
sram_add_entry(0, 4, 684, 4, 128'h40300000000000000000000ea98);
sram_add_entry(0, 4, 688, 4, 128'h403000000000000000000008e43);
sram_add_entry(0, 4, 692, 4, 128'h403000000000000000000002164);
sram_add_entry(0, 4, 696, 4, 128'h403000000000000000000003319);
sram_add_entry(0, 4, 700, 4, 128'h40300000000000000000000a7d4);
sram_add_entry(0, 4, 704, 4, 128'h4030000000000000000000032a8);
sram_add_entry(0, 4, 708, 4, 128'h40300000000000000000000e83b);
sram_add_entry(0, 4, 712, 4, 128'h403000000000000000000001fb9);
sram_add_entry(0, 4, 716, 4, 128'h4030000000000000000000097e4);
sram_add_entry(0, 4, 720, 4, 128'h40300000000000000000000c832);
sram_add_entry(0, 4, 724, 4, 128'h403000000000000000000004045);
sram_add_entry(0, 4, 728, 4, 128'h403000000000000000000002e4b);
sram_add_entry(0, 4, 732, 4, 128'h403000000000000000000005001);
sram_add_entry(0, 4, 736, 4, 128'h4030000000000000000000089f4);
sram_add_entry(0, 4, 740, 4, 128'h403000000000000000000004f20);
sram_add_entry(0, 4, 744, 4, 128'h40300000000000000000000718d);
sram_add_entry(0, 4, 748, 4, 128'h40300000000000000000000ec81);
sram_add_entry(0, 4, 752, 4, 128'h40300000000000000000000eff2);
sram_add_entry(0, 4, 756, 4, 128'h4030000000000000000000032f9);
sram_add_entry(0, 4, 760, 4, 128'h40300000000000000000000df51);
sram_add_entry(0, 4, 764, 4, 128'h40300000000000000000000aebe);
sram_add_entry(0, 4, 768, 4, 128'h403000000000000000000001952);
sram_add_entry(0, 4, 772, 4, 128'h40300000000000000000000989a);
sram_add_entry(0, 4, 776, 4, 128'h403000000000000000000004d90);
sram_add_entry(0, 4, 780, 4, 128'h40300000000000000000000cda6);
sram_add_entry(0, 4, 784, 4, 128'h4030000000000000000000011cf);
sram_add_entry(0, 4, 788, 4, 128'h4030000000000000000000046d5);
sram_add_entry(0, 4, 792, 4, 128'h40300000000000000000000cdeb);
sram_add_entry(0, 4, 796, 4, 128'h4030000000000000000000060b3);
sram_add_entry(0, 4, 800, 4, 128'h40300000000000000000000e8cc);
sram_add_entry(0, 4, 804, 4, 128'h4030000000000000000000099ed);
sram_add_entry(0, 4, 808, 4, 128'h40300000000000000000000c9aa);
sram_add_entry(0, 4, 812, 4, 128'h40300000000000000000000a401);
sram_add_entry(0, 4, 816, 4, 128'h40300000000000000000000a4a0);
sram_add_entry(0, 4, 820, 4, 128'h403000000000000000000009821);
sram_add_entry(0, 4, 824, 4, 128'h40300000000000000000000e330);
sram_add_entry(0, 4, 828, 4, 128'h403000000000000000000005327);
sram_add_entry(0, 4, 832, 4, 128'h40300000000000000000000085c);
sram_add_entry(0, 4, 836, 4, 128'h40300000000000000000000f8ea);
sram_add_entry(0, 4, 840, 4, 128'h40300000000000000000000243d);
sram_add_entry(0, 4, 844, 4, 128'h4030000000000000000000067f8);
sram_add_entry(0, 4, 848, 4, 128'h4030000000000000000000055bf);
sram_add_entry(0, 4, 852, 4, 128'h40300000000000000000000731b);
sram_add_entry(0, 4, 856, 4, 128'h4030000000000000000000080fd);
sram_add_entry(0, 4, 860, 4, 128'h40300000000000000000000af4c);
sram_add_entry(0, 4, 864, 4, 128'h403000000000000000000004a57);
sram_add_entry(0, 4, 868, 4, 128'h40300000000000000000000414d);
sram_add_entry(0, 4, 872, 4, 128'h403000000000000000000005dd0);
sram_add_entry(0, 4, 876, 4, 128'h403000000000000000000007720);
sram_add_entry(0, 4, 880, 4, 128'h40300000000000000000000378c);
sram_add_entry(0, 4, 884, 4, 128'h40300000000000000000000c49c);
sram_add_entry(0, 4, 888, 4, 128'h4030000000000000000000097f4);
sram_add_entry(0, 4, 892, 4, 128'h403000000000000000000007335);
sram_add_entry(0, 4, 896, 4, 128'h40300000000000000000000130f);
sram_add_entry(0, 4, 900, 4, 128'h403000000000000000000009dc0);
sram_add_entry(0, 4, 904, 4, 128'h40300000000000000000000f760);
sram_add_entry(0, 4, 908, 4, 128'h403000000000000000000001800);
sram_add_entry(0, 4, 912, 4, 128'h4030000000000000000000040fe);
sram_add_entry(0, 4, 916, 4, 128'h40300000000000000000000698d);
sram_add_entry(0, 4, 920, 4, 128'h40300000000000000000000ac63);
sram_add_entry(0, 4, 924, 4, 128'h403000000000000000000000cb0);
sram_add_entry(0, 4, 928, 4, 128'h40300000000000000000000a762);
sram_add_entry(0, 4, 932, 4, 128'h40300000000000000000000c7e3);
sram_add_entry(0, 4, 936, 4, 128'h403000000000000000000007950);
sram_add_entry(0, 4, 940, 4, 128'h40300000000000000000000393f);
sram_add_entry(0, 4, 944, 4, 128'h40300000000000000000000b5a0);
sram_add_entry(0, 4, 948, 4, 128'h40300000000000000000000a992);
sram_add_entry(0, 4, 952, 4, 128'h403000000000000000000009d82);
sram_add_entry(0, 4, 956, 4, 128'h403000000000000000000004659);
sram_add_entry(0, 4, 960, 4, 128'h4030000000000000000000099f3);
sram_add_entry(0, 4, 964, 4, 128'h4030000000000000000000031f6);
sram_add_entry(0, 4, 968, 4, 128'h403000000000000000000004389);
sram_add_entry(0, 4, 972, 4, 128'h403000000000000000000009fbe);
sram_add_entry(0, 4, 976, 4, 128'h403000000000000000000001fa1);
sram_add_entry(0, 4, 980, 4, 128'h403000000000000000000004eb0);
sram_add_entry(0, 4, 984, 4, 128'h40300000000000000000000af41);
sram_add_entry(0, 4, 988, 4, 128'h403000000000000000000008b0d);
sram_add_entry(0, 4, 992, 4, 128'h40300000000000000000000b721);
sram_add_entry(0, 4, 996, 4, 128'h40300000000000000000000b055);
sram_add_entry(0, 4, 1000, 4, 128'h40300000000000000000000a3fa);
sram_add_entry(0, 4, 1004, 4, 128'h40300000000000000000000f530);
sram_add_entry(0, 4, 1008, 4, 128'h4030000000000000000000040ec);
sram_add_entry(0, 4, 1012, 4, 128'h40300000000000000000000bf82);
sram_add_entry(0, 4, 1016, 4, 128'h403000000000000000000002613);
sram_add_entry(0, 4, 1020, 4, 128'h403000000000000000000007010);
sram_add_entry(0, 4, 1024, 4, 128'h40300000000000000000000c20c);
sram_add_entry(0, 4, 1028, 4, 128'h40300000000000000000000b5a2);
sram_add_entry(0, 4, 1032, 4, 128'h4030000000000000000000007d6);
sram_add_entry(0, 4, 1036, 4, 128'h403000000000000000000008c9b);
sram_add_entry(0, 4, 1040, 4, 128'h403000000000000000000002cb2);
sram_add_entry(0, 4, 1044, 4, 128'h40300000000000000000000ac1b);
sram_add_entry(0, 4, 1048, 4, 128'h40300000000000000000000c493);
sram_add_entry(0, 4, 1052, 4, 128'h403000000000000000000002fc6);
sram_add_entry(0, 4, 1056, 4, 128'h40300000000000000000000a2b9);
sram_add_entry(0, 4, 1060, 4, 128'h40300000000000000000000f03a);
sram_add_entry(0, 4, 1064, 4, 128'h40300000000000000000000628c);
sram_add_entry(0, 4, 1068, 4, 128'h403000000000000000000008a4f);
sram_add_entry(0, 4, 1072, 4, 128'h40300000000000000000000f6ce);
sram_add_entry(0, 4, 1076, 4, 128'h4030000000000000000000094f6);
sram_add_entry(0, 4, 1080, 4, 128'h403000000000000000000005ff0);
sram_add_entry(0, 4, 1084, 4, 128'h40300000000000000000000dd7f);
sram_add_entry(0, 4, 1088, 4, 128'h40300000000000000000000e12f);
sram_add_entry(0, 4, 1092, 4, 128'h40300000000000000000000773e);
sram_add_entry(0, 4, 1096, 4, 128'h40300000000000000000000add4);
sram_add_entry(0, 4, 1100, 4, 128'h40300000000000000000000bc61);
sram_add_entry(0, 4, 1104, 4, 128'h40300000000000000000000bce1);
sram_add_entry(0, 4, 1108, 4, 128'h403000000000000000000007c3d);
sram_add_entry(0, 4, 1112, 4, 128'h40300000000000000000000cbb3);
sram_add_entry(0, 4, 1116, 4, 128'h4030000000000000000000047e1);
sram_add_entry(0, 4, 1120, 4, 128'h4030000000000000000000054ac);
sram_add_entry(0, 4, 1124, 4, 128'h403000000000000000000000d99);
sram_add_entry(0, 4, 1128, 4, 128'h40300000000000000000000337c);
sram_add_entry(0, 4, 1132, 4, 128'h4030000000000000000000070b8);
sram_add_entry(0, 4, 1136, 4, 128'h40300000000000000000000732e);
sram_add_entry(0, 4, 1140, 4, 128'h403000000000000000000006d44);
sram_add_entry(0, 4, 1144, 4, 128'h403000000000000000000005f66);
sram_add_entry(0, 4, 1148, 4, 128'h40300000000000000000000cead);
sram_add_entry(0, 4, 1152, 4, 128'h4030000000000000000000035a7);
sram_add_entry(0, 4, 1156, 4, 128'h4030000000000000000000036bd);
sram_add_entry(0, 4, 1160, 4, 128'h403000000000000000000009924);
sram_add_entry(0, 4, 1164, 4, 128'h403000000000000000000009e17);
sram_add_entry(0, 4, 1168, 4, 128'h40300000000000000000000c72a);
sram_add_entry(0, 4, 1172, 4, 128'h403000000000000000000004ee3);
sram_add_entry(0, 4, 1176, 4, 128'h4030000000000000000000005e7);
sram_add_entry(0, 4, 1180, 4, 128'h40300000000000000000000b1e7);
sram_add_entry(0, 4, 1184, 4, 128'h403000000000000000000005cac);
sram_add_entry(0, 4, 1188, 4, 128'h403000000000000000000007c98);
sram_add_entry(0, 4, 1192, 4, 128'h40300000000000000000000f24a);
sram_add_entry(0, 4, 1196, 4, 128'h403000000000000000000009017);
sram_add_entry(0, 4, 1200, 4, 128'h403000000000000000000000a86);
sram_add_entry(0, 4, 1204, 4, 128'h4030000000000000000000015c7);
sram_add_entry(0, 4, 1208, 4, 128'h403000000000000000000006c3d);
sram_add_entry(0, 4, 1212, 4, 128'h40300000000000000000000501e);
sram_add_entry(0, 4, 1216, 4, 128'h4030000000000000000000010c9);
sram_add_entry(0, 4, 1220, 4, 128'h403000000000000000000005862);
sram_add_entry(0, 4, 1224, 4, 128'h40300000000000000000000028e);
sram_add_entry(0, 4, 1228, 4, 128'h40300000000000000000000c850);
sram_add_entry(0, 4, 1232, 4, 128'h40300000000000000000000af6c);
sram_add_entry(0, 4, 1236, 4, 128'h4030000000000000000000090d3);
sram_add_entry(0, 4, 1240, 4, 128'h40300000000000000000000b6b1);
sram_add_entry(0, 4, 1244, 4, 128'h403000000000000000000005e8d);
sram_add_entry(0, 4, 1248, 4, 128'h403000000000000000000005855);
sram_add_entry(0, 4, 1252, 4, 128'h403000000000000000000006c01);
sram_add_entry(0, 4, 1256, 4, 128'h40300000000000000000000dcb4);
sram_add_entry(0, 4, 1260, 4, 128'h40300000000000000000000c207);
sram_add_entry(0, 4, 1264, 4, 128'h40300000000000000000000f4c7);
sram_add_entry(0, 4, 1268, 4, 128'h40300000000000000000000c655);
sram_add_entry(0, 4, 1272, 4, 128'h403000000000000000000005a6a);
sram_add_entry(0, 4, 1276, 4, 128'h40300000000000000000000fdf1);
sram_add_entry(0, 4, 1280, 4, 128'h40300000000000000000000762c);
sram_add_entry(0, 4, 1284, 4, 128'h403000000000000000000003342);
sram_add_entry(0, 4, 1288, 4, 128'h40300000000000000000000a47d);
sram_add_entry(0, 4, 1292, 4, 128'h40300000000000000000000049d);
sram_add_entry(0, 4, 1296, 4, 128'h403000000000000000000004c88);
sram_add_entry(0, 4, 1300, 4, 128'h40300000000000000000000b9a2);
sram_add_entry(0, 4, 1304, 4, 128'h40300000000000000000000605b);
sram_add_entry(0, 4, 1308, 4, 128'h403000000000000000000001b57);
sram_add_entry(0, 4, 1312, 4, 128'h403000000000000000000002d7c);
sram_add_entry(0, 4, 1316, 4, 128'h40300000000000000000000598d);
sram_add_entry(0, 4, 1320, 4, 128'h40300000000000000000000bad0);
sram_add_entry(0, 4, 1324, 4, 128'h403000000000000000000002246);
sram_add_entry(0, 4, 1328, 4, 128'h40300000000000000000000a559);
sram_add_entry(0, 4, 1332, 4, 128'h40300000000000000000000e9bd);
sram_add_entry(0, 4, 1336, 4, 128'h40300000000000000000000ba7c);
sram_add_entry(0, 4, 1340, 4, 128'h40300000000000000000000bf4e);
sram_add_entry(0, 4, 1344, 4, 128'h40300000000000000000000505a);
sram_add_entry(0, 4, 1348, 4, 128'h403000000000000000000007213);
sram_add_entry(0, 4, 1352, 4, 128'h403000000000000000000007e6d);
sram_add_entry(0, 4, 1356, 4, 128'h40300000000000000000000676e);
sram_add_entry(0, 4, 1360, 4, 128'h40300000000000000000000191f);
sram_add_entry(0, 4, 1364, 4, 128'h403000000000000000000003181);
sram_add_entry(0, 4, 1368, 4, 128'h4030000000000000000000017ab);
sram_add_entry(0, 4, 1372, 4, 128'h403000000000000000000003075);
sram_add_entry(0, 4, 1376, 4, 128'h40300000000000000000000afc7);
sram_add_entry(0, 4, 1380, 4, 128'h40300000000000000000000cde1);
sram_add_entry(0, 4, 1384, 4, 128'h403000000000000000000004ffc);
sram_add_entry(0, 4, 1388, 4, 128'h40300000000000000000000dc23);
sram_add_entry(0, 4, 1392, 4, 128'h403000000000000000000000d21);
sram_add_entry(0, 4, 1396, 4, 128'h403000000000000000000006432);
sram_add_entry(0, 4, 1400, 4, 128'h40300000000000000000000925a);
sram_add_entry(0, 4, 1404, 4, 128'h40300000000000000000000c72e);
sram_add_entry(0, 4, 1408, 4, 128'h4030000000000000000000059d9);
sram_add_entry(0, 4, 1412, 4, 128'h403000000000000000000007e41);
sram_add_entry(0, 4, 1416, 4, 128'h40300000000000000000000e51e);
sram_add_entry(0, 4, 1420, 4, 128'h403000000000000000000002182);
sram_add_entry(0, 4, 1424, 4, 128'h4030000000000000000000085fd);
sram_add_entry(0, 4, 1428, 4, 128'h40300000000000000000000ff81);
sram_add_entry(0, 4, 1432, 4, 128'h40300000000000000000000abc8);
sram_add_entry(0, 4, 1436, 4, 128'h403000000000000000000000933);
sram_add_entry(0, 4, 1440, 4, 128'h40300000000000000000000075b);
sram_add_entry(0, 4, 1444, 4, 128'h40300000000000000000000e194);
sram_add_entry(0, 4, 1448, 4, 128'h40300000000000000000000a000);
sram_add_entry(0, 4, 1452, 4, 128'h4030000000000000000000075d7);
sram_add_entry(0, 4, 1456, 4, 128'h403000000000000000000002796);
sram_add_entry(0, 4, 1460, 4, 128'h40300000000000000000000e2de);
sram_add_entry(0, 4, 1464, 4, 128'h40300000000000000000000fb48);
sram_add_entry(0, 4, 1468, 4, 128'h403000000000000000000006be4);
sram_add_entry(0, 4, 1472, 4, 128'h403000000000000000000000a2f);
sram_add_entry(0, 4, 1476, 4, 128'h403000000000000000000008b4f);
sram_add_entry(0, 4, 1480, 4, 128'h40300000000000000000000f592);
sram_add_entry(0, 4, 1484, 4, 128'h403000000000000000000002cc7);
sram_add_entry(0, 4, 1488, 4, 128'h40300000000000000000000b053);
sram_add_entry(0, 4, 1492, 4, 128'h40300000000000000000000a982);
sram_add_entry(0, 4, 1496, 4, 128'h40300000000000000000000f7f5);
sram_add_entry(0, 4, 1500, 4, 128'h40300000000000000000000abff);
sram_add_entry(0, 4, 1504, 4, 128'h40300000000000000000000c5a1);
sram_add_entry(0, 4, 1508, 4, 128'h40300000000000000000000c504);
sram_add_entry(0, 4, 1512, 4, 128'h40300000000000000000000260b);
sram_add_entry(0, 4, 1516, 4, 128'h40300000000000000000000ecef);
sram_add_entry(0, 4, 1520, 4, 128'h403000000000000000000001548);
sram_add_entry(0, 4, 1524, 4, 128'h4030000000000000000000063f7);
sram_add_entry(0, 4, 1528, 4, 128'h40300000000000000000000097c);
sram_add_entry(0, 4, 1532, 4, 128'h40300000000000000000000492e);
sram_add_entry(0, 4, 1536, 4, 128'h403000000000000000000007d91);
sram_add_entry(0, 4, 1540, 4, 128'h403000000000000000000005e33);
sram_add_entry(0, 4, 1544, 4, 128'h4030000000000000000000020ff);
sram_add_entry(0, 4, 1548, 4, 128'h403000000000000000000002d2b);
sram_add_entry(0, 4, 1552, 4, 128'h403000000000000000000004faf);
sram_add_entry(0, 4, 1556, 4, 128'h403000000000000000000009fc0);
sram_add_entry(0, 4, 1560, 4, 128'h403000000000000000000007df6);
sram_add_entry(0, 4, 1564, 4, 128'h403000000000000000000008145);
sram_add_entry(0, 4, 1568, 4, 128'h40300000000000000000000d8dc);
sram_add_entry(0, 4, 1572, 4, 128'h403000000000000000000008ccb);
sram_add_entry(0, 4, 1576, 4, 128'h40300000000000000000000a74c);
sram_add_entry(0, 4, 1580, 4, 128'h40300000000000000000000d54d);
sram_add_entry(0, 4, 1584, 4, 128'h4030000000000000000000057ec);
sram_add_entry(0, 4, 1588, 4, 128'h40300000000000000000000d895);
sram_add_entry(0, 4, 1592, 4, 128'h403000000000000000000004a8a);
sram_add_entry(0, 4, 1596, 4, 128'h40300000000000000000000aad5);
sram_add_entry(0, 4, 1600, 4, 128'h403000000000000000000002dc8);
sram_add_entry(0, 4, 1604, 4, 128'h40300000000000000000000d305);
sram_add_entry(0, 4, 1608, 4, 128'h40300000000000000000000f654);
sram_add_entry(0, 4, 1612, 4, 128'h403000000000000000000007cef);
sram_add_entry(0, 4, 1616, 4, 128'h40300000000000000000000fdcd);
sram_add_entry(0, 4, 1620, 4, 128'h403000000000000000000009c53);
sram_add_entry(0, 4, 1624, 4, 128'h4030000000000000000000056bf);
sram_add_entry(0, 4, 1628, 4, 128'h40300000000000000000000df03);
sram_add_entry(0, 4, 1632, 4, 128'h403000000000000000000008eb7);
sram_add_entry(0, 4, 1636, 4, 128'h4030000000000000000000027c4);
sram_add_entry(0, 4, 1640, 4, 128'h403000000000000000000006ae4);
sram_add_entry(0, 4, 1644, 4, 128'h403000000000000000000008beb);
sram_add_entry(0, 4, 1648, 4, 128'h403000000000000000000006ac7);
sram_add_entry(0, 4, 1652, 4, 128'h40300000000000000000000c8ce);
sram_add_entry(0, 4, 1656, 4, 128'h403000000000000000000000f6f);
sram_add_entry(0, 4, 1660, 4, 128'h40300000000000000000000c185);
sram_add_entry(0, 4, 1664, 4, 128'h403000000000000000000008ecb);
sram_add_entry(0, 4, 1668, 4, 128'h40300000000000000000000c088);
sram_add_entry(0, 4, 1672, 4, 128'h40300000000000000000000fb13);
sram_add_entry(0, 4, 1676, 4, 128'h403000000000000000000008323);
sram_add_entry(0, 4, 1680, 4, 128'h4030000000000000000000004be);
sram_add_entry(0, 4, 1684, 4, 128'h40300000000000000000000d5d8);
sram_add_entry(0, 4, 1688, 4, 128'h40300000000000000000000f5e5);
sram_add_entry(0, 4, 1692, 4, 128'h40300000000000000000000e858);
sram_add_entry(0, 4, 1696, 4, 128'h40300000000000000000000ec83);
sram_add_entry(0, 4, 1700, 4, 128'h403000000000000000000004b57);
sram_add_entry(0, 4, 1704, 4, 128'h403000000000000000000007510);
sram_add_entry(0, 4, 1708, 4, 128'h403000000000000000000007e0c);
sram_add_entry(0, 4, 1712, 4, 128'h40300000000000000000000afdd);
sram_add_entry(0, 4, 1716, 4, 128'h40300000000000000000000eea0);
sram_add_entry(0, 4, 1720, 4, 128'h40300000000000000000000dc6b);
sram_add_entry(0, 4, 1724, 4, 128'h40300000000000000000000dc6d);
sram_add_entry(0, 4, 1728, 4, 128'h40300000000000000000000f267);
sram_add_entry(0, 4, 1732, 4, 128'h40300000000000000000000cc96);
sram_add_entry(0, 4, 1736, 4, 128'h403000000000000000000006e0e);
sram_add_entry(0, 4, 1740, 4, 128'h40300000000000000000000adf2);
sram_add_entry(0, 4, 1744, 4, 128'h4030000000000000000000022cf);
sram_add_entry(0, 4, 1748, 4, 128'h40300000000000000000000efe3);
sram_add_entry(0, 4, 1752, 4, 128'h40300000000000000000000327f);
sram_add_entry(0, 4, 1756, 4, 128'h40300000000000000000000c1cd);
sram_add_entry(0, 4, 1760, 4, 128'h4030000000000000000000087d7);
sram_add_entry(0, 4, 1764, 4, 128'h4030000000000000000000052ae);
sram_add_entry(0, 4, 1768, 4, 128'h40300000000000000000000522d);
sram_add_entry(0, 4, 1772, 4, 128'h4030000000000000000000023e9);
sram_add_entry(0, 4, 1776, 4, 128'h403000000000000000000009f00);
sram_add_entry(0, 4, 1780, 4, 128'h403000000000000000000004222);
sram_add_entry(0, 4, 1784, 4, 128'h40300000000000000000000c826);
sram_add_entry(0, 4, 1788, 4, 128'h403000000000000000000005c33);
sram_add_entry(0, 4, 1792, 4, 128'h4030000000000000000000025c2);
sram_add_entry(0, 4, 1796, 4, 128'h40300000000000000000000c4f6);
sram_add_entry(0, 4, 1800, 4, 128'h40300000000000000000000f947);
sram_add_entry(0, 4, 1804, 4, 128'h4030000000000000000000075e1);
sram_add_entry(0, 4, 1808, 4, 128'h403000000000000000000004b59);
sram_add_entry(0, 4, 1812, 4, 128'h40300000000000000000000cc5d);
sram_add_entry(0, 4, 1816, 4, 128'h40300000000000000000000ec89);
sram_add_entry(0, 4, 1820, 4, 128'h40300000000000000000000ac8e);
sram_add_entry(0, 4, 1824, 4, 128'h403000000000000000000009306);
sram_add_entry(0, 4, 1828, 4, 128'h40300000000000000000000b015);
sram_add_entry(0, 4, 1832, 4, 128'h403000000000000000000009893);
sram_add_entry(0, 4, 1836, 4, 128'h40300000000000000000000a323);
sram_add_entry(0, 4, 1840, 4, 128'h403000000000000000000002482);
sram_add_entry(0, 4, 1844, 4, 128'h4030000000000000000000073ba);
sram_add_entry(0, 4, 1848, 4, 128'h403000000000000000000008241);
sram_add_entry(0, 4, 1852, 4, 128'h4030000000000000000000002c7);
sram_add_entry(0, 4, 1856, 4, 128'h403000000000000000000003d42);
sram_add_entry(0, 4, 1860, 4, 128'h4030000000000000000000009b8);
sram_add_entry(0, 4, 1864, 4, 128'h403000000000000000000006583);
sram_add_entry(0, 4, 1868, 4, 128'h40300000000000000000000e989);
sram_add_entry(0, 4, 1872, 4, 128'h4030000000000000000000077b8);
sram_add_entry(0, 4, 1876, 4, 128'h40300000000000000000000372f);
sram_add_entry(0, 4, 1880, 4, 128'h40300000000000000000000ef75);
sram_add_entry(0, 4, 1884, 4, 128'h40300000000000000000000e2a0);
sram_add_entry(0, 4, 1888, 4, 128'h40300000000000000000000f84a);
sram_add_entry(0, 4, 1892, 4, 128'h40300000000000000000000e2f5);
sram_add_entry(0, 4, 1896, 4, 128'h40300000000000000000000ca43);
sram_add_entry(0, 4, 1900, 4, 128'h40300000000000000000000b85f);
sram_add_entry(0, 4, 1904, 4, 128'h40300000000000000000000b9fd);
sram_add_entry(0, 4, 1908, 4, 128'h40300000000000000000000730d);
sram_add_entry(0, 4, 1912, 4, 128'h40300000000000000000000bd98);
sram_add_entry(0, 4, 1916, 4, 128'h403000000000000000000007046);
sram_add_entry(0, 4, 1920, 4, 128'h40300000000000000000000c7f0);
sram_add_entry(0, 4, 1924, 4, 128'h403000000000000000000007b74);
sram_add_entry(0, 4, 1928, 4, 128'h40300000000000000000000117f);
sram_add_entry(0, 4, 1932, 4, 128'h40300000000000000000000a024);
sram_add_entry(0, 4, 1936, 4, 128'h40300000000000000000000b6cc);
sram_add_entry(0, 4, 1940, 4, 128'h403000000000000000000005a3f);
sram_add_entry(0, 4, 1944, 4, 128'h40300000000000000000000bf61);
sram_add_entry(0, 4, 1948, 4, 128'h40300000000000000000000c96b);
sram_add_entry(0, 4, 1952, 4, 128'h40300000000000000000000c476);
sram_add_entry(0, 4, 1956, 4, 128'h40300000000000000000000c029);
sram_add_entry(0, 4, 1960, 4, 128'h40300000000000000000000446f);
sram_add_entry(0, 4, 1964, 4, 128'h40300000000000000000000c986);
sram_add_entry(0, 4, 1968, 4, 128'h403000000000000000000008bf2);
sram_add_entry(0, 4, 1972, 4, 128'h40300000000000000000000190b);
sram_add_entry(0, 4, 1976, 4, 128'h403000000000000000000002afd);
sram_add_entry(0, 4, 1980, 4, 128'h403000000000000000000009aad);
sram_add_entry(0, 4, 1984, 4, 128'h40300000000000000000000e797);
sram_add_entry(0, 4, 1988, 4, 128'h40300000000000000000000c09a);
sram_add_entry(0, 4, 1992, 4, 128'h40300000000000000000000671f);
sram_add_entry(0, 4, 1996, 4, 128'h403000000000000000000004c2c);
sram_add_entry(0, 4, 2000, 4, 128'h403000000000000000000003ef1);
sram_add_entry(0, 4, 2004, 4, 128'h40300000000000000000000c600);
sram_add_entry(0, 4, 2008, 4, 128'h403000000000000000000006ce5);
sram_add_entry(0, 4, 2012, 4, 128'h403000000000000000000001228);
sram_add_entry(0, 4, 2016, 4, 128'h40300000000000000000000e80e);
sram_add_entry(0, 4, 2020, 4, 128'h403000000000000000000008dd7);
sram_add_entry(0, 4, 2024, 4, 128'h40300000000000000000000d9ff);
sram_add_entry(0, 4, 2028, 4, 128'h403000000000000000000009114);
sram_add_entry(0, 4, 2032, 4, 128'h40300000000000000000000fffd);
sram_add_entry(0, 4, 2036, 4, 128'h40300000000000000000000fec1);
sram_add_entry(0, 4, 2040, 4, 128'h40300000000000000000000157a);
sram_add_entry(0, 4, 2044, 4, 128'h403000000000000000000008698);
sram_add_entry(0, 4, 2048, 4, 128'h4030000000000000000000064dd);
sram_add_entry(0, 4, 2052, 4, 128'h403000000000000000000006c7b);
sram_add_entry(0, 4, 2056, 4, 128'h40300000000000000000000d6f6);
sram_add_entry(0, 4, 2060, 4, 128'h40300000000000000000000d74e);
sram_add_entry(0, 4, 2064, 4, 128'h40300000000000000000000d5ca);
sram_add_entry(0, 4, 2068, 4, 128'h403000000000000000000007199);
sram_add_entry(0, 4, 2072, 4, 128'h403000000000000000000005167);
sram_add_entry(0, 4, 2076, 4, 128'h403000000000000000000002b74);
sram_add_entry(0, 4, 2080, 4, 128'h40300000000000000000000418b);
sram_add_entry(0, 4, 2084, 4, 128'h403000000000000000000004e9a);
sram_add_entry(0, 4, 2088, 4, 128'h403000000000000000000008692);
sram_add_entry(0, 4, 2092, 4, 128'h40300000000000000000000c6e0);
sram_add_entry(0, 4, 2096, 4, 128'h403000000000000000000001f44);
sram_add_entry(0, 4, 2100, 4, 128'h4030000000000000000000075a0);
sram_add_entry(0, 4, 2104, 4, 128'h403000000000000000000003793);
sram_add_entry(0, 4, 2108, 4, 128'h403000000000000000000006365);
sram_add_entry(0, 4, 2112, 4, 128'h40300000000000000000000ee99);
sram_add_entry(0, 4, 2116, 4, 128'h403000000000000000000000ac5);
sram_add_entry(0, 4, 2120, 4, 128'h403000000000000000000006b09);
sram_add_entry(0, 4, 2124, 4, 128'h4030000000000000000000054d0);
sram_add_entry(0, 4, 2128, 4, 128'h40300000000000000000000b98d);
sram_add_entry(0, 4, 2132, 4, 128'h40300000000000000000000d586);
sram_add_entry(0, 4, 2136, 4, 128'h403000000000000000000004cc3);
sram_add_entry(0, 4, 2140, 4, 128'h40300000000000000000000c26c);
sram_add_entry(0, 4, 2144, 4, 128'h40300000000000000000000f681);
sram_add_entry(0, 4, 2148, 4, 128'h40300000000000000000000f0c9);
sram_add_entry(0, 4, 2152, 4, 128'h40300000000000000000000be02);
sram_add_entry(0, 4, 2156, 4, 128'h403000000000000000000005eb8);
sram_add_entry(0, 4, 2160, 4, 128'h403000000000000000000004c1e);
sram_add_entry(0, 4, 2164, 4, 128'h40300000000000000000000c52a);
sram_add_entry(0, 4, 2168, 4, 128'h40300000000000000000000093c);
sram_add_entry(0, 4, 2172, 4, 128'h40300000000000000000000d07f);
sram_add_entry(0, 4, 2176, 4, 128'h40300000000000000000000d767);
sram_add_entry(0, 4, 2180, 4, 128'h4030000000000000000000029db);
sram_add_entry(0, 4, 2184, 4, 128'h403000000000000000000002546);
sram_add_entry(0, 4, 2188, 4, 128'h4030000000000000000000012d9);
sram_add_entry(0, 4, 2192, 4, 128'h40300000000000000000000ff67);
sram_add_entry(0, 4, 2196, 4, 128'h40300000000000000000000da73);
sram_add_entry(0, 4, 2200, 4, 128'h403000000000000000000000b6d);
sram_add_entry(0, 4, 2204, 4, 128'h40300000000000000000000f5b5);
sram_add_entry(0, 4, 2208, 4, 128'h4030000000000000000000006e7);
sram_add_entry(0, 4, 2212, 4, 128'h40300000000000000000000d236);
sram_add_entry(0, 4, 2216, 4, 128'h40300000000000000000000b505);
sram_add_entry(0, 4, 2220, 4, 128'h403000000000000000000007813);
sram_add_entry(0, 4, 2224, 4, 128'h40300000000000000000000199a);
sram_add_entry(0, 4, 2228, 4, 128'h403000000000000000000001e9d);
sram_add_entry(0, 4, 2232, 4, 128'h403000000000000000000008438);
sram_add_entry(0, 4, 2236, 4, 128'h40300000000000000000000853c);
sram_add_entry(0, 4, 2240, 4, 128'h40300000000000000000000fa90);
sram_add_entry(0, 4, 2244, 4, 128'h4030000000000000000000091d3);
sram_add_entry(0, 4, 2248, 4, 128'h403000000000000000000009871);
sram_add_entry(0, 4, 2252, 4, 128'h40300000000000000000000f155);
sram_add_entry(0, 4, 2256, 4, 128'h403000000000000000000000ec3);
sram_add_entry(0, 4, 2260, 4, 128'h403000000000000000000000240);
sram_add_entry(0, 4, 2264, 4, 128'h40300000000000000000000c7bf);
sram_add_entry(0, 4, 2268, 4, 128'h403000000000000000000003579);
sram_add_entry(0, 4, 2272, 4, 128'h403000000000000000000006f16);
sram_add_entry(0, 4, 2276, 4, 128'h403000000000000000000002fbd);
sram_add_entry(0, 4, 2280, 4, 128'h40300000000000000000000376f);
sram_add_entry(0, 4, 2284, 4, 128'h403000000000000000000008129);
sram_add_entry(0, 4, 2288, 4, 128'h40300000000000000000000cb9c);
sram_add_entry(0, 4, 2292, 4, 128'h403000000000000000000008b5a);
sram_add_entry(0, 4, 2296, 4, 128'h40300000000000000000000c137);
sram_add_entry(0, 4, 2300, 4, 128'h4030000000000000000000016b5);
sram_add_entry(0, 4, 2304, 4, 128'h403000000000000000000009006);
sram_add_entry(0, 4, 2308, 4, 128'h4030000000000000000000024fd);
sram_add_entry(0, 4, 2312, 4, 128'h4030000000000000000000038c7);
sram_add_entry(0, 4, 2316, 4, 128'h40300000000000000000000f065);
sram_add_entry(0, 4, 2320, 4, 128'h40300000000000000000000d149);
sram_add_entry(0, 4, 2324, 4, 128'h40300000000000000000000f573);
sram_add_entry(0, 4, 2328, 4, 128'h40300000000000000000000a7e5);
sram_add_entry(0, 4, 2332, 4, 128'h40300000000000000000000c110);
sram_add_entry(0, 4, 2336, 4, 128'h403000000000000000000006859);
sram_add_entry(0, 4, 2340, 4, 128'h4030000000000000000000066bb);
sram_add_entry(0, 4, 2344, 4, 128'h403000000000000000000006dc2);
sram_add_entry(0, 4, 2348, 4, 128'h40300000000000000000000fce5);
sram_add_entry(0, 4, 2352, 4, 128'h4030000000000000000000089f3);
sram_add_entry(0, 4, 2356, 4, 128'h40300000000000000000000188f);
sram_add_entry(0, 4, 2360, 4, 128'h403000000000000000000000c76);
sram_add_entry(0, 4, 2364, 4, 128'h403000000000000000000000d66);
sram_add_entry(0, 4, 2368, 4, 128'h403000000000000000000008a86);
sram_add_entry(0, 4, 2372, 4, 128'h403000000000000000000002056);
sram_add_entry(0, 4, 2376, 4, 128'h40300000000000000000000c598);
sram_add_entry(0, 4, 2380, 4, 128'h403000000000000000000001cb6);
sram_add_entry(0, 4, 2384, 4, 128'h4030000000000000000000079c6);
sram_add_entry(0, 4, 2388, 4, 128'h403000000000000000000007621);
sram_add_entry(0, 4, 2392, 4, 128'h40300000000000000000000bd5d);
sram_add_entry(0, 4, 2396, 4, 128'h4030000000000000000000080e8);
sram_add_entry(0, 4, 2400, 4, 128'h40300000000000000000000581f);
sram_add_entry(0, 4, 2404, 4, 128'h40300000000000000000000c915);
sram_add_entry(0, 4, 2408, 4, 128'h403000000000000000000001142);
sram_add_entry(0, 4, 2412, 4, 128'h4030000000000000000000039df);
sram_add_entry(0, 4, 2416, 4, 128'h4030000000000000000000055cc);
sram_add_entry(0, 4, 2420, 4, 128'h40300000000000000000000f2a1);
sram_add_entry(0, 4, 2424, 4, 128'h40300000000000000000000fa13);
sram_add_entry(0, 4, 2428, 4, 128'h4030000000000000000000004c4);
sram_add_entry(0, 4, 2432, 4, 128'h40300000000000000000000aa67);
sram_add_entry(0, 4, 2436, 4, 128'h40300000000000000000000187a);
sram_add_entry(0, 4, 2440, 4, 128'h403000000000000000000008437);
sram_add_entry(0, 4, 2444, 4, 128'h403000000000000000000000faf);
sram_add_entry(0, 4, 2448, 4, 128'h4030000000000000000000010bb);
sram_add_entry(0, 4, 2452, 4, 128'h40300000000000000000000c03c);
sram_add_entry(0, 4, 2456, 4, 128'h40300000000000000000000a17d);
sram_add_entry(0, 4, 2460, 4, 128'h40300000000000000000000a172);
sram_add_entry(0, 4, 2464, 4, 128'h4030000000000000000000036c5);
sram_add_entry(0, 4, 2468, 4, 128'h40300000000000000000000344d);
sram_add_entry(0, 4, 2472, 4, 128'h403000000000000000000004e82);
sram_add_entry(0, 4, 2476, 4, 128'h40300000000000000000000e473);
sram_add_entry(0, 4, 2480, 4, 128'h403000000000000000000004bfd);
sram_add_entry(0, 4, 2484, 4, 128'h40300000000000000000000d436);
sram_add_entry(0, 4, 2488, 4, 128'h4030000000000000000000033a7);
sram_add_entry(0, 4, 2492, 4, 128'h40300000000000000000000e4bf);
sram_add_entry(0, 4, 2496, 4, 128'h403000000000000000000004c20);
sram_add_entry(0, 4, 2500, 4, 128'h40300000000000000000000c7cc);
sram_add_entry(0, 4, 2504, 4, 128'h403000000000000000000002ff0);
sram_add_entry(0, 4, 2508, 4, 128'h4030000000000000000000033c8);
sram_add_entry(0, 4, 2512, 4, 128'h4030000000000000000000040c4);
sram_add_entry(0, 4, 2516, 4, 128'h4030000000000000000000064a9);
sram_add_entry(0, 4, 2520, 4, 128'h40300000000000000000000078d);
sram_add_entry(0, 4, 2524, 4, 128'h40300000000000000000000a2d3);
sram_add_entry(0, 4, 2528, 4, 128'h403000000000000000000003326);
sram_add_entry(0, 4, 2532, 4, 128'h40300000000000000000000dbf9);
sram_add_entry(0, 4, 2536, 4, 128'h40300000000000000000000907a);
sram_add_entry(0, 4, 2540, 4, 128'h40300000000000000000000e187);
sram_add_entry(0, 4, 2544, 4, 128'h403000000000000000000001c66);
sram_add_entry(0, 4, 2548, 4, 128'h40300000000000000000000f67e);
sram_add_entry(0, 4, 2552, 4, 128'h403000000000000000000004aa1);
sram_add_entry(0, 4, 2556, 4, 128'h40300000000000000000000fd6b);
sram_add_entry(0, 4, 2560, 4, 128'h40300000000000000000000b65b);
sram_add_entry(0, 4, 2564, 4, 128'h4030000000000000000000050f8);
sram_add_entry(0, 4, 2568, 4, 128'h40300000000000000000000ee03);
sram_add_entry(0, 4, 2572, 4, 128'h40300000000000000000000bf2d);
sram_add_entry(0, 4, 2576, 4, 128'h403000000000000000000005809);
sram_add_entry(0, 4, 2580, 4, 128'h40300000000000000000000e9a7);
sram_add_entry(0, 4, 2584, 4, 128'h40300000000000000000000f3f3);
sram_add_entry(0, 4, 2588, 4, 128'h403000000000000000000008ce2);
sram_add_entry(0, 4, 2592, 4, 128'h40300000000000000000000c953);
sram_add_entry(0, 4, 2596, 4, 128'h403000000000000000000000b0d);
sram_add_entry(0, 4, 2600, 4, 128'h40300000000000000000000623b);
sram_add_entry(0, 4, 2604, 4, 128'h40300000000000000000000a57a);
sram_add_entry(0, 4, 2608, 4, 128'h40300000000000000000000bbfd);
sram_add_entry(0, 4, 2612, 4, 128'h403000000000000000000000cd5);
sram_add_entry(0, 4, 2616, 4, 128'h4030000000000000000000007d9);
sram_add_entry(0, 4, 2620, 4, 128'h40300000000000000000000d5b7);
sram_add_entry(0, 4, 2624, 4, 128'h40300000000000000000000c765);
sram_add_entry(0, 4, 2628, 4, 128'h40300000000000000000000af71);
sram_add_entry(0, 4, 2632, 4, 128'h40300000000000000000000e0e2);
sram_add_entry(0, 4, 2636, 4, 128'h40300000000000000000000eab4);
sram_add_entry(0, 4, 2640, 4, 128'h40300000000000000000000b006);
sram_add_entry(0, 4, 2644, 4, 128'h40300000000000000000000a268);
sram_add_entry(0, 4, 2648, 4, 128'h403000000000000000000002e18);
sram_add_entry(0, 4, 2652, 4, 128'h403000000000000000000008f7d);
sram_add_entry(0, 4, 2656, 4, 128'h40300000000000000000000b733);
sram_add_entry(0, 4, 2660, 4, 128'h403000000000000000000007454);
sram_add_entry(0, 4, 2664, 4, 128'h403000000000000000000000651);
sram_add_entry(0, 4, 2668, 4, 128'h4030000000000000000000021c7);
sram_add_entry(0, 4, 2672, 4, 128'h40300000000000000000000f615);
sram_add_entry(0, 4, 2676, 4, 128'h40300000000000000000000d932);
sram_add_entry(0, 4, 2680, 4, 128'h40300000000000000000000dc24);
sram_add_entry(0, 4, 2684, 4, 128'h403000000000000000000006b3b);
sram_add_entry(0, 4, 2688, 4, 128'h40300000000000000000000a575);
sram_add_entry(0, 4, 2692, 4, 128'h403000000000000000000007f07);
sram_add_entry(0, 4, 2696, 4, 128'h40300000000000000000000bb77);
sram_add_entry(0, 4, 2700, 4, 128'h403000000000000000000004308);
sram_add_entry(0, 4, 2704, 4, 128'h40300000000000000000000901d);
sram_add_entry(0, 4, 2708, 4, 128'h403000000000000000000002f04);
sram_add_entry(0, 4, 2712, 4, 128'h403000000000000000000000672);
sram_add_entry(0, 4, 2716, 4, 128'h403000000000000000000004440);
sram_add_entry(0, 4, 2720, 4, 128'h403000000000000000000000222);
sram_add_entry(0, 4, 2724, 4, 128'h40300000000000000000000208f);
sram_add_entry(0, 4, 2728, 4, 128'h40300000000000000000000b0a7);
sram_add_entry(0, 4, 2732, 4, 128'h403000000000000000000001a32);
sram_add_entry(0, 4, 2736, 4, 128'h40300000000000000000000b3cd);
sram_add_entry(0, 4, 2740, 4, 128'h40300000000000000000000cef3);
sram_add_entry(0, 4, 2744, 4, 128'h403000000000000000000005f33);
sram_add_entry(0, 4, 2748, 4, 128'h403000000000000000000005003);
sram_add_entry(0, 4, 2752, 4, 128'h403000000000000000000002cb3);
sram_add_entry(0, 4, 2756, 4, 128'h40300000000000000000000f670);
sram_add_entry(0, 4, 2760, 4, 128'h40300000000000000000000b8be);
sram_add_entry(0, 4, 2764, 4, 128'h40300000000000000000000254b);
sram_add_entry(0, 4, 2768, 4, 128'h40300000000000000000000b525);
sram_add_entry(0, 4, 2772, 4, 128'h403000000000000000000009a07);
sram_add_entry(0, 4, 2776, 4, 128'h40300000000000000000000af14);
sram_add_entry(0, 4, 2780, 4, 128'h40300000000000000000000759e);
sram_add_entry(0, 4, 2784, 4, 128'h40300000000000000000000d9b5);
sram_add_entry(0, 4, 2788, 4, 128'h403000000000000000000002612);
sram_add_entry(0, 4, 2792, 4, 128'h40300000000000000000000e49c);
sram_add_entry(0, 4, 2796, 4, 128'h40300000000000000000000fc4a);
sram_add_entry(0, 4, 2800, 4, 128'h40300000000000000000000d6fd);
