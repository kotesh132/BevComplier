initial
begin
sos_loop[0].somModel.tcam_data[1][0][0]=80'h00000000000000000000;
sos_loop[0].somModel.tcam_mask[1][0][0]=80'hffffffffffffffffffff;
sos_loop[0].somModel.tcam_data[1][1][0]=80'h000000009b2571c7073c;
sos_loop[0].somModel.tcam_mask[1][1][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][2][0]=80'h00000000ede35ed4bae4;
sos_loop[0].somModel.tcam_mask[1][2][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][3][0]=80'h00000000d835b1486b13;
sos_loop[0].somModel.tcam_mask[1][3][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][4][0]=80'h00000000be3dd6d14071;
sos_loop[0].somModel.tcam_mask[1][4][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][5][0]=80'h0000000088e0f6aa248a;
sos_loop[0].somModel.tcam_mask[1][5][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][6][0]=80'h00000000f3012b605570;
sos_loop[0].somModel.tcam_mask[1][6][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][7][0]=80'h00000000e16202381133;
sos_loop[0].somModel.tcam_mask[1][7][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][8][0]=80'h00000000f16aa927fb4a;
sos_loop[0].somModel.tcam_mask[1][8][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][9][0]=80'h00000000458011f44fab;
sos_loop[0].somModel.tcam_mask[1][9][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][10][0]=80'h000000006b5603b74017;
sos_loop[0].somModel.tcam_mask[1][10][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][11][0]=80'h000000009867863b5169;
sos_loop[0].somModel.tcam_mask[1][11][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][12][0]=80'h000000007d563611e661;
sos_loop[0].somModel.tcam_mask[1][12][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][13][0]=80'h000000009a388934f048;
sos_loop[0].somModel.tcam_mask[1][13][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][14][0]=80'h00000000e7d208135786;
sos_loop[0].somModel.tcam_mask[1][14][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][15][0]=80'h000000001d236be012e4;
sos_loop[0].somModel.tcam_mask[1][15][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][16][0]=80'h0000000004816ad6457a;
sos_loop[0].somModel.tcam_mask[1][16][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[1][17][0]=80'h00000000b7fcfacfa875;
sos_loop[0].somModel.tcam_mask[1][17][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][18][0]=80'h00000000acdaf0aca7c6;
sos_loop[0].somModel.tcam_mask[1][18][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][19][0]=80'h00000000272061475aea;
sos_loop[0].somModel.tcam_mask[1][19][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][20][0]=80'h00000000ed5c1ad98d27;
sos_loop[0].somModel.tcam_mask[1][20][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][21][0]=80'h0000000005137add3842;
sos_loop[0].somModel.tcam_mask[1][21][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[1][22][0]=80'h0000000077c13eb8f0bc;
sos_loop[0].somModel.tcam_mask[1][22][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][23][0]=80'h0000000064dec849f297;
sos_loop[0].somModel.tcam_mask[1][23][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][24][0]=80'h0000000052815aaa0e76;
sos_loop[0].somModel.tcam_mask[1][24][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][25][0]=80'h0000000036c627639625;
sos_loop[0].somModel.tcam_mask[1][25][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][26][0]=80'h00000000adfa0e35ab63;
sos_loop[0].somModel.tcam_mask[1][26][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][27][0]=80'h00000000de873f211f1b;
sos_loop[0].somModel.tcam_mask[1][27][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][28][0]=80'h000000007c056a29eb06;
sos_loop[0].somModel.tcam_mask[1][28][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][29][0]=80'h00000000b17370ad5889;
sos_loop[0].somModel.tcam_mask[1][29][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][30][0]=80'h000000003c16a3b80a77;
sos_loop[0].somModel.tcam_mask[1][30][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][31][0]=80'h00000000fdc75e2fe46f;
sos_loop[0].somModel.tcam_mask[1][31][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][32][0]=80'h00000000b514aca9a7ea;
sos_loop[0].somModel.tcam_mask[1][32][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][33][0]=80'h00000000ff4fc0b5dd4f;
sos_loop[0].somModel.tcam_mask[1][33][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][34][0]=80'h000000004fa3edb32414;
sos_loop[0].somModel.tcam_mask[1][34][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][35][0]=80'h00000000a7a0a91df8ba;
sos_loop[0].somModel.tcam_mask[1][35][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][36][0]=80'h00000000f1dccb540bd9;
sos_loop[0].somModel.tcam_mask[1][36][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][37][0]=80'h00000000db32f0046c0d;
sos_loop[0].somModel.tcam_mask[1][37][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][38][0]=80'h000000005be7f8e59bc2;
sos_loop[0].somModel.tcam_mask[1][38][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][39][0]=80'h0000000056ae936d2b74;
sos_loop[0].somModel.tcam_mask[1][39][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][40][0]=80'h0000000021237dd3755f;
sos_loop[0].somModel.tcam_mask[1][40][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][41][0]=80'h00000000a6839f79036b;
sos_loop[0].somModel.tcam_mask[1][41][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][42][0]=80'h0000000005e54e001a27;
sos_loop[0].somModel.tcam_mask[1][42][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[1][43][0]=80'h000000002dfc19bbb79a;
sos_loop[0].somModel.tcam_mask[1][43][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][44][0]=80'h000000007da11a068ee0;
sos_loop[0].somModel.tcam_mask[1][44][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][45][0]=80'h000000007b392b497f6e;
sos_loop[0].somModel.tcam_mask[1][45][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][46][0]=80'h000000006c0398426174;
sos_loop[0].somModel.tcam_mask[1][46][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][47][0]=80'h000000007b724903d7a9;
sos_loop[0].somModel.tcam_mask[1][47][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][48][0]=80'h000000007e2e109e6271;
sos_loop[0].somModel.tcam_mask[1][48][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][49][0]=80'h0000000070b0857e229f;
sos_loop[0].somModel.tcam_mask[1][49][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][50][0]=80'h00000000276af0ce7d95;
sos_loop[0].somModel.tcam_mask[1][50][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][51][0]=80'h00000000977c2662d661;
sos_loop[0].somModel.tcam_mask[1][51][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][52][0]=80'h000000006c110a6ebb5c;
sos_loop[0].somModel.tcam_mask[1][52][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][53][0]=80'h000000007100f4f63c98;
sos_loop[0].somModel.tcam_mask[1][53][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][54][0]=80'h000000000dee6b07e350;
sos_loop[0].somModel.tcam_mask[1][54][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][55][0]=80'h0000000073f1bab9b30b;
sos_loop[0].somModel.tcam_mask[1][55][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][56][0]=80'h0000000045a7a7cd7c56;
sos_loop[0].somModel.tcam_mask[1][56][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][57][0]=80'h000000005c2982129594;
sos_loop[0].somModel.tcam_mask[1][57][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][58][0]=80'h0000000024f31697e85b;
sos_loop[0].somModel.tcam_mask[1][58][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][59][0]=80'h000000001217e5938719;
sos_loop[0].somModel.tcam_mask[1][59][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][60][0]=80'h00000000d7165d2854bd;
sos_loop[0].somModel.tcam_mask[1][60][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][61][0]=80'h00000000a943cd77303b;
sos_loop[0].somModel.tcam_mask[1][61][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][62][0]=80'h00000000eb90c7477f53;
sos_loop[0].somModel.tcam_mask[1][62][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][63][0]=80'h00000000445c3e0895fe;
sos_loop[0].somModel.tcam_mask[1][63][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][64][0]=80'h00000000b312060a0eef;
sos_loop[0].somModel.tcam_mask[1][64][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][65][0]=80'h00000000cc66a816d743;
sos_loop[0].somModel.tcam_mask[1][65][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][66][0]=80'h00000000b3497a7141e9;
sos_loop[0].somModel.tcam_mask[1][66][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][67][0]=80'h00000000822765751942;
sos_loop[0].somModel.tcam_mask[1][67][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][68][0]=80'h00000000199ff6767d07;
sos_loop[0].somModel.tcam_mask[1][68][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][69][0]=80'h00000000d15a97c2415f;
sos_loop[0].somModel.tcam_mask[1][69][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][70][0]=80'h00000000e029b33bdf0c;
sos_loop[0].somModel.tcam_mask[1][70][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][71][0]=80'h00000000516f120d3a96;
sos_loop[0].somModel.tcam_mask[1][71][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][72][0]=80'h000000004e9aec95e85c;
sos_loop[0].somModel.tcam_mask[1][72][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][73][0]=80'h00000000d172c141c22a;
sos_loop[0].somModel.tcam_mask[1][73][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][74][0]=80'h0000000073147f2a5ee0;
sos_loop[0].somModel.tcam_mask[1][74][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][75][0]=80'h00000000fbb8275391e0;
sos_loop[0].somModel.tcam_mask[1][75][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][76][0]=80'h0000000065fdd1b8aab4;
sos_loop[0].somModel.tcam_mask[1][76][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][77][0]=80'h00000000f1874d4b4c76;
sos_loop[0].somModel.tcam_mask[1][77][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][78][0]=80'h000000006cd16dcc4a33;
sos_loop[0].somModel.tcam_mask[1][78][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][79][0]=80'h00000000d96441dc2078;
sos_loop[0].somModel.tcam_mask[1][79][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][80][0]=80'h00000000c319811fd277;
sos_loop[0].somModel.tcam_mask[1][80][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][81][0]=80'h000000008a0471dd6d11;
sos_loop[0].somModel.tcam_mask[1][81][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][82][0]=80'h00000000f394863f8076;
sos_loop[0].somModel.tcam_mask[1][82][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][83][0]=80'h000000005b121b7039e5;
sos_loop[0].somModel.tcam_mask[1][83][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][84][0]=80'h00000000eafeaba615dc;
sos_loop[0].somModel.tcam_mask[1][84][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][85][0]=80'h00000000c10aef68e81f;
sos_loop[0].somModel.tcam_mask[1][85][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][86][0]=80'h00000000b4285b984022;
sos_loop[0].somModel.tcam_mask[1][86][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][87][0]=80'h000000008264ffadb985;
sos_loop[0].somModel.tcam_mask[1][87][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][88][0]=80'h000000000a5638ebc9ea;
sos_loop[0].somModel.tcam_mask[1][88][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][89][0]=80'h00000000c025ca05681b;
sos_loop[0].somModel.tcam_mask[1][89][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][90][0]=80'h0000000069fc597ace55;
sos_loop[0].somModel.tcam_mask[1][90][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][91][0]=80'h0000000092d13ceb35ee;
sos_loop[0].somModel.tcam_mask[1][91][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][92][0]=80'h00000000d92c798e2da4;
sos_loop[0].somModel.tcam_mask[1][92][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][93][0]=80'h00000000ef44bbde26b8;
sos_loop[0].somModel.tcam_mask[1][93][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][94][0]=80'h000000004a7bde16a1b0;
sos_loop[0].somModel.tcam_mask[1][94][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][95][0]=80'h000000009cef75742606;
sos_loop[0].somModel.tcam_mask[1][95][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][96][0]=80'h00000000bc689291a89e;
sos_loop[0].somModel.tcam_mask[1][96][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][97][0]=80'h00000000ecad85584eac;
sos_loop[0].somModel.tcam_mask[1][97][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][98][0]=80'h000000002596ab0bd4ef;
sos_loop[0].somModel.tcam_mask[1][98][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][99][0]=80'h00000000afb0bcd5f28c;
sos_loop[0].somModel.tcam_mask[1][99][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][100][0]=80'h00000000588ea274f953;
sos_loop[0].somModel.tcam_mask[1][100][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][101][0]=80'h00000000a7391453de54;
sos_loop[0].somModel.tcam_mask[1][101][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][102][0]=80'h00000000fdbcbd10e033;
sos_loop[0].somModel.tcam_mask[1][102][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][103][0]=80'h00000000719cfa2767c3;
sos_loop[0].somModel.tcam_mask[1][103][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][104][0]=80'h00000000a3ef35e42c33;
sos_loop[0].somModel.tcam_mask[1][104][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][105][0]=80'h00000000c4c69a60a71a;
sos_loop[0].somModel.tcam_mask[1][105][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][106][0]=80'h000000003a3a7b0a793b;
sos_loop[0].somModel.tcam_mask[1][106][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][107][0]=80'h00000000cfa4b3cac05c;
sos_loop[0].somModel.tcam_mask[1][107][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][108][0]=80'h000000005599e50df8a9;
sos_loop[0].somModel.tcam_mask[1][108][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][109][0]=80'h000000003a0f6debddd0;
sos_loop[0].somModel.tcam_mask[1][109][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][110][0]=80'h000000009f11ab78573a;
sos_loop[0].somModel.tcam_mask[1][110][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][111][0]=80'h00000000d608068e6320;
sos_loop[0].somModel.tcam_mask[1][111][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][112][0]=80'h00000000d862045cf75f;
sos_loop[0].somModel.tcam_mask[1][112][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][113][0]=80'h000000006cae027bae23;
sos_loop[0].somModel.tcam_mask[1][113][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][114][0]=80'h00000000e2a567e44491;
sos_loop[0].somModel.tcam_mask[1][114][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][115][0]=80'h0000000072c9f8b64ee2;
sos_loop[0].somModel.tcam_mask[1][115][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][116][0]=80'h00000000408440fab4cd;
sos_loop[0].somModel.tcam_mask[1][116][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][117][0]=80'h000000004309898b60f3;
sos_loop[0].somModel.tcam_mask[1][117][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][118][0]=80'h00000000115a7eb75e3a;
sos_loop[0].somModel.tcam_mask[1][118][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][119][0]=80'h0000000037178729e67f;
sos_loop[0].somModel.tcam_mask[1][119][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][120][0]=80'h00000000fb424524db25;
sos_loop[0].somModel.tcam_mask[1][120][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][121][0]=80'h00000000361984d7eb12;
sos_loop[0].somModel.tcam_mask[1][121][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][122][0]=80'h00000000927e86180bf1;
sos_loop[0].somModel.tcam_mask[1][122][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][123][0]=80'h000000006a2879654a57;
sos_loop[0].somModel.tcam_mask[1][123][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][124][0]=80'h00000000641b343f80f4;
sos_loop[0].somModel.tcam_mask[1][124][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][125][0]=80'h0000000093991f1d7362;
sos_loop[0].somModel.tcam_mask[1][125][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][126][0]=80'h0000000015e87559900d;
sos_loop[0].somModel.tcam_mask[1][126][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][127][0]=80'h000000005d613c992175;
sos_loop[0].somModel.tcam_mask[1][127][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][128][0]=80'h00000000899161eca21b;
sos_loop[0].somModel.tcam_mask[1][128][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][129][0]=80'h000000004a353e6fdb65;
sos_loop[0].somModel.tcam_mask[1][129][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][130][0]=80'h000000006d2289d6b1b5;
sos_loop[0].somModel.tcam_mask[1][130][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][131][0]=80'h0000000063d6892f4cbd;
sos_loop[0].somModel.tcam_mask[1][131][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][132][0]=80'h000000000ec516e56e38;
sos_loop[0].somModel.tcam_mask[1][132][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][133][0]=80'h00000000f6d75e867538;
sos_loop[0].somModel.tcam_mask[1][133][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][134][0]=80'h00000000f8103fe52fca;
sos_loop[0].somModel.tcam_mask[1][134][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][135][0]=80'h000000003721758992ed;
sos_loop[0].somModel.tcam_mask[1][135][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][136][0]=80'h00000000c7a4b46ded9a;
sos_loop[0].somModel.tcam_mask[1][136][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][137][0]=80'h000000008261693eedaf;
sos_loop[0].somModel.tcam_mask[1][137][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][138][0]=80'h000000003a70bd4ccb71;
sos_loop[0].somModel.tcam_mask[1][138][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][139][0]=80'h00000000dc3e4883a653;
sos_loop[0].somModel.tcam_mask[1][139][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][140][0]=80'h000000006bb7508ac2dc;
sos_loop[0].somModel.tcam_mask[1][140][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][141][0]=80'h00000000873638a207ca;
sos_loop[0].somModel.tcam_mask[1][141][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][142][0]=80'h0000000004732c91bc5c;
sos_loop[0].somModel.tcam_mask[1][142][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[1][143][0]=80'h000000003fd9b4c00a99;
sos_loop[0].somModel.tcam_mask[1][143][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][144][0]=80'h00000000859aa75fc399;
sos_loop[0].somModel.tcam_mask[1][144][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][145][0]=80'h0000000078ba5e9eee08;
sos_loop[0].somModel.tcam_mask[1][145][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][146][0]=80'h0000000000dbd3b819af;
sos_loop[0].somModel.tcam_mask[1][146][0]=80'hffffffffff0000000000;
sos_loop[0].somModel.tcam_data[1][147][0]=80'h00000000080957200a77;
sos_loop[0].somModel.tcam_mask[1][147][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][148][0]=80'h00000000ad807c006574;
sos_loop[0].somModel.tcam_mask[1][148][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][149][0]=80'h00000000b25671eb1928;
sos_loop[0].somModel.tcam_mask[1][149][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][150][0]=80'h00000000cd733d038007;
sos_loop[0].somModel.tcam_mask[1][150][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][151][0]=80'h000000005a808481d4f8;
sos_loop[0].somModel.tcam_mask[1][151][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][152][0]=80'h00000000e5270474bc3d;
sos_loop[0].somModel.tcam_mask[1][152][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][153][0]=80'h0000000043c133e30238;
sos_loop[0].somModel.tcam_mask[1][153][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][154][0]=80'h00000000da06327c0fb6;
sos_loop[0].somModel.tcam_mask[1][154][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][155][0]=80'h00000000f44aa55e8d5b;
sos_loop[0].somModel.tcam_mask[1][155][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][156][0]=80'h00000000d108767b16e2;
sos_loop[0].somModel.tcam_mask[1][156][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][157][0]=80'h0000000045b722c61027;
sos_loop[0].somModel.tcam_mask[1][157][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][158][0]=80'h00000000a633db8c75b8;
sos_loop[0].somModel.tcam_mask[1][158][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][159][0]=80'h00000000f2d4b44fd6dc;
sos_loop[0].somModel.tcam_mask[1][159][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][160][0]=80'h00000000affaa97c08bb;
sos_loop[0].somModel.tcam_mask[1][160][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][161][0]=80'h000000003db1f6e4e6a5;
sos_loop[0].somModel.tcam_mask[1][161][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][162][0]=80'h00000000cc8499d91df3;
sos_loop[0].somModel.tcam_mask[1][162][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][163][0]=80'h00000000bde381c08689;
sos_loop[0].somModel.tcam_mask[1][163][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][164][0]=80'h000000004903fd0700cd;
sos_loop[0].somModel.tcam_mask[1][164][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][165][0]=80'h000000001af8bbb7c7be;
sos_loop[0].somModel.tcam_mask[1][165][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][166][0]=80'h00000000d7cd2a4ee374;
sos_loop[0].somModel.tcam_mask[1][166][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][167][0]=80'h00000000648e675ea632;
sos_loop[0].somModel.tcam_mask[1][167][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][168][0]=80'h0000000002ab6d3cad9b;
sos_loop[0].somModel.tcam_mask[1][168][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[1][169][0]=80'h000000005f26b6f13520;
sos_loop[0].somModel.tcam_mask[1][169][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][170][0]=80'h00000000a96772107053;
sos_loop[0].somModel.tcam_mask[1][170][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][171][0]=80'h00000000fd5134dc543a;
sos_loop[0].somModel.tcam_mask[1][171][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][172][0]=80'h00000000f9e15e388cda;
sos_loop[0].somModel.tcam_mask[1][172][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][173][0]=80'h0000000037ad0dd04d1b;
sos_loop[0].somModel.tcam_mask[1][173][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][174][0]=80'h0000000024ed9e62765c;
sos_loop[0].somModel.tcam_mask[1][174][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][175][0]=80'h00000000deaa2a8e2c76;
sos_loop[0].somModel.tcam_mask[1][175][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][176][0]=80'h000000009afd8ccdf0d3;
sos_loop[0].somModel.tcam_mask[1][176][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][177][0]=80'h00000000dfba92cc34c0;
sos_loop[0].somModel.tcam_mask[1][177][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][178][0]=80'h000000001d1b77568814;
sos_loop[0].somModel.tcam_mask[1][178][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][179][0]=80'h00000000c138abed4b17;
sos_loop[0].somModel.tcam_mask[1][179][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][180][0]=80'h0000000038fe88806ab3;
sos_loop[0].somModel.tcam_mask[1][180][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][181][0]=80'h00000000f4a91c35928f;
sos_loop[0].somModel.tcam_mask[1][181][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][182][0]=80'h0000000053d53e8897d5;
sos_loop[0].somModel.tcam_mask[1][182][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][183][0]=80'h0000000091213c03913d;
sos_loop[0].somModel.tcam_mask[1][183][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][184][0]=80'h0000000039beec93c1a6;
sos_loop[0].somModel.tcam_mask[1][184][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][185][0]=80'h00000000b842fcc92642;
sos_loop[0].somModel.tcam_mask[1][185][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][186][0]=80'h000000005350a885c6e9;
sos_loop[0].somModel.tcam_mask[1][186][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][187][0]=80'h000000003a60895d3611;
sos_loop[0].somModel.tcam_mask[1][187][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][188][0]=80'h000000003958522de12b;
sos_loop[0].somModel.tcam_mask[1][188][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][189][0]=80'h000000008379dd2f10a6;
sos_loop[0].somModel.tcam_mask[1][189][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][190][0]=80'h00000000719a6a66e65a;
sos_loop[0].somModel.tcam_mask[1][190][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][191][0]=80'h00000000151b0bccc299;
sos_loop[0].somModel.tcam_mask[1][191][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][192][0]=80'h0000000060a3a0ebb851;
sos_loop[0].somModel.tcam_mask[1][192][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][193][0]=80'h00000000ceeb751d2978;
sos_loop[0].somModel.tcam_mask[1][193][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][194][0]=80'h000000006799c24bb3b7;
sos_loop[0].somModel.tcam_mask[1][194][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][195][0]=80'h0000000056badc0db157;
sos_loop[0].somModel.tcam_mask[1][195][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][196][0]=80'h000000004feefc3e7730;
sos_loop[0].somModel.tcam_mask[1][196][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][197][0]=80'h00000000d3f5a6c1574e;
sos_loop[0].somModel.tcam_mask[1][197][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][198][0]=80'h00000000b6364f27da3b;
sos_loop[0].somModel.tcam_mask[1][198][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][199][0]=80'h00000000df1f0128cbbd;
sos_loop[0].somModel.tcam_mask[1][199][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][200][0]=80'h0000000009cd060e84aa;
sos_loop[0].somModel.tcam_mask[1][200][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][201][0]=80'h000000008373ac34c47f;
sos_loop[0].somModel.tcam_mask[1][201][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][202][0]=80'h000000001e386f8b863d;
sos_loop[0].somModel.tcam_mask[1][202][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][203][0]=80'h000000005ba2afce95f3;
sos_loop[0].somModel.tcam_mask[1][203][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][204][0]=80'h000000004e2599a1897a;
sos_loop[0].somModel.tcam_mask[1][204][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][205][0]=80'h00000000f5479d3b77c5;
sos_loop[0].somModel.tcam_mask[1][205][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][206][0]=80'h00000000abbe127976b8;
sos_loop[0].somModel.tcam_mask[1][206][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][207][0]=80'h00000000da3b98564520;
sos_loop[0].somModel.tcam_mask[1][207][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][208][0]=80'h000000005ac0acc44533;
sos_loop[0].somModel.tcam_mask[1][208][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][209][0]=80'h00000000ddd77ea80899;
sos_loop[0].somModel.tcam_mask[1][209][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][210][0]=80'h000000005ab30dbacc5d;
sos_loop[0].somModel.tcam_mask[1][210][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][211][0]=80'h00000000342220f18625;
sos_loop[0].somModel.tcam_mask[1][211][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][212][0]=80'h000000002a04827b867b;
sos_loop[0].somModel.tcam_mask[1][212][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][213][0]=80'h00000000541f28ab2585;
sos_loop[0].somModel.tcam_mask[1][213][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][214][0]=80'h00000000283b331b6fc3;
sos_loop[0].somModel.tcam_mask[1][214][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][215][0]=80'h000000006f3ac91b9a16;
sos_loop[0].somModel.tcam_mask[1][215][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][216][0]=80'h0000000041fd7e0e3811;
sos_loop[0].somModel.tcam_mask[1][216][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][217][0]=80'h0000000058966af35810;
sos_loop[0].somModel.tcam_mask[1][217][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][218][0]=80'h00000000e9cafeeb8643;
sos_loop[0].somModel.tcam_mask[1][218][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][219][0]=80'h00000000b3e98f6adfb5;
sos_loop[0].somModel.tcam_mask[1][219][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][220][0]=80'h00000000739e76de29f1;
sos_loop[0].somModel.tcam_mask[1][220][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][221][0]=80'h000000002a304169ea35;
sos_loop[0].somModel.tcam_mask[1][221][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][222][0]=80'h000000008151be21591a;
sos_loop[0].somModel.tcam_mask[1][222][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][223][0]=80'h000000001225f462349c;
sos_loop[0].somModel.tcam_mask[1][223][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][224][0]=80'h000000002719c0ef3496;
sos_loop[0].somModel.tcam_mask[1][224][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][225][0]=80'h0000000054fb7f3c0cef;
sos_loop[0].somModel.tcam_mask[1][225][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][226][0]=80'h00000000fef0454047a7;
sos_loop[0].somModel.tcam_mask[1][226][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][227][0]=80'h00000000b4d08228d18c;
sos_loop[0].somModel.tcam_mask[1][227][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][228][0]=80'h00000000a167559cde76;
sos_loop[0].somModel.tcam_mask[1][228][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][229][0]=80'h0000000093813f42c579;
sos_loop[0].somModel.tcam_mask[1][229][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][230][0]=80'h000000008510d813599c;
sos_loop[0].somModel.tcam_mask[1][230][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][231][0]=80'h00000000d983360209d9;
sos_loop[0].somModel.tcam_mask[1][231][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][232][0]=80'h000000009b211b4fc467;
sos_loop[0].somModel.tcam_mask[1][232][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][233][0]=80'h000000002330c01b4962;
sos_loop[0].somModel.tcam_mask[1][233][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][234][0]=80'h00000000844df8e1f63b;
sos_loop[0].somModel.tcam_mask[1][234][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][235][0]=80'h00000000c041ca14cdca;
sos_loop[0].somModel.tcam_mask[1][235][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][236][0]=80'h00000000daae12e7d039;
sos_loop[0].somModel.tcam_mask[1][236][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][237][0]=80'h000000007036cba3dc70;
sos_loop[0].somModel.tcam_mask[1][237][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][238][0]=80'h00000000f19f6d156eb4;
sos_loop[0].somModel.tcam_mask[1][238][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][239][0]=80'h0000000089fcfce01525;
sos_loop[0].somModel.tcam_mask[1][239][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][240][0]=80'h000000001fad9639ae38;
sos_loop[0].somModel.tcam_mask[1][240][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][241][0]=80'h0000000059882292a37d;
sos_loop[0].somModel.tcam_mask[1][241][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][242][0]=80'h00000000d1c038664adc;
sos_loop[0].somModel.tcam_mask[1][242][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][243][0]=80'h0000000050d6e9dd8cb9;
sos_loop[0].somModel.tcam_mask[1][243][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][244][0]=80'h0000000068165950944c;
sos_loop[0].somModel.tcam_mask[1][244][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][245][0]=80'h00000000b1b417cc4d0d;
sos_loop[0].somModel.tcam_mask[1][245][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][246][0]=80'h00000000673c0c16111e;
sos_loop[0].somModel.tcam_mask[1][246][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][247][0]=80'h000000009282fc16753b;
sos_loop[0].somModel.tcam_mask[1][247][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][248][0]=80'h000000000465552830d4;
sos_loop[0].somModel.tcam_mask[1][248][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[1][249][0]=80'h00000000a237c12459ce;
sos_loop[0].somModel.tcam_mask[1][249][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][250][0]=80'h000000003fbff4f63ebe;
sos_loop[0].somModel.tcam_mask[1][250][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][251][0]=80'h0000000083622bea46ac;
sos_loop[0].somModel.tcam_mask[1][251][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][252][0]=80'h00000000ace489475745;
sos_loop[0].somModel.tcam_mask[1][252][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][253][0]=80'h000000001b62f58d5c3b;
sos_loop[0].somModel.tcam_mask[1][253][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][254][0]=80'h000000003d317dd9a17e;
sos_loop[0].somModel.tcam_mask[1][254][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][255][0]=80'h000000009b4487a8ad15;
sos_loop[0].somModel.tcam_mask[1][255][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][256][0]=80'h000000001eb8f0ced706;
sos_loop[0].somModel.tcam_mask[1][256][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][257][0]=80'h0000000023df27639b89;
sos_loop[0].somModel.tcam_mask[1][257][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][258][0]=80'h000000009e02d67f2c49;
sos_loop[0].somModel.tcam_mask[1][258][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][259][0]=80'h000000002f03370d25d5;
sos_loop[0].somModel.tcam_mask[1][259][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][260][0]=80'h0000000023c475b331f3;
sos_loop[0].somModel.tcam_mask[1][260][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][261][0]=80'h000000000298cf5b269e;
sos_loop[0].somModel.tcam_mask[1][261][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[1][262][0]=80'h00000000e8d802a6eec6;
sos_loop[0].somModel.tcam_mask[1][262][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][263][0]=80'h00000000b112320fcf2c;
sos_loop[0].somModel.tcam_mask[1][263][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][264][0]=80'h000000001e8b12608817;
sos_loop[0].somModel.tcam_mask[1][264][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][265][0]=80'h0000000070b74d52680c;
sos_loop[0].somModel.tcam_mask[1][265][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][266][0]=80'h000000009385b9ebc706;
sos_loop[0].somModel.tcam_mask[1][266][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][267][0]=80'h00000000c5ddaac7946a;
sos_loop[0].somModel.tcam_mask[1][267][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][268][0]=80'h00000000d71073217127;
sos_loop[0].somModel.tcam_mask[1][268][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][269][0]=80'h00000000d100d643c643;
sos_loop[0].somModel.tcam_mask[1][269][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][270][0]=80'h00000000f69ca57a9df0;
sos_loop[0].somModel.tcam_mask[1][270][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][271][0]=80'h00000000ff6881bbfec2;
sos_loop[0].somModel.tcam_mask[1][271][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][272][0]=80'h00000000f2823e7062c6;
sos_loop[0].somModel.tcam_mask[1][272][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][273][0]=80'h0000000061e0198f5ae3;
sos_loop[0].somModel.tcam_mask[1][273][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][274][0]=80'h000000002693612b76f7;
sos_loop[0].somModel.tcam_mask[1][274][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][275][0]=80'h000000009e4433b3d0ed;
sos_loop[0].somModel.tcam_mask[1][275][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][276][0]=80'h000000001aa909a924ce;
sos_loop[0].somModel.tcam_mask[1][276][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][277][0]=80'h000000000529bf4b7234;
sos_loop[0].somModel.tcam_mask[1][277][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[1][278][0]=80'h0000000071c5876f6f41;
sos_loop[0].somModel.tcam_mask[1][278][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][279][0]=80'h000000004840ebc670dd;
sos_loop[0].somModel.tcam_mask[1][279][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][280][0]=80'h00000000e8a44e161d3a;
sos_loop[0].somModel.tcam_mask[1][280][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][281][0]=80'h0000000045616bb46ded;
sos_loop[0].somModel.tcam_mask[1][281][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][282][0]=80'h0000000052dcbdb0812e;
sos_loop[0].somModel.tcam_mask[1][282][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][283][0]=80'h0000000074514d0e52f1;
sos_loop[0].somModel.tcam_mask[1][283][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][284][0]=80'h0000000095635f45a99d;
sos_loop[0].somModel.tcam_mask[1][284][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][285][0]=80'h000000007ec8277acb2c;
sos_loop[0].somModel.tcam_mask[1][285][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][286][0]=80'h000000000df530f8507d;
sos_loop[0].somModel.tcam_mask[1][286][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][287][0]=80'h0000000076c5dc4ff347;
sos_loop[0].somModel.tcam_mask[1][287][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][288][0]=80'h00000000da63394fdb26;
sos_loop[0].somModel.tcam_mask[1][288][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][289][0]=80'h00000000df60cec8ddc2;
sos_loop[0].somModel.tcam_mask[1][289][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][290][0]=80'h00000000777e53ca6502;
sos_loop[0].somModel.tcam_mask[1][290][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][291][0]=80'h00000000fa9ef6faf654;
sos_loop[0].somModel.tcam_mask[1][291][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][292][0]=80'h00000000e2fa7ff677c6;
sos_loop[0].somModel.tcam_mask[1][292][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][293][0]=80'h000000001a6d4480a388;
sos_loop[0].somModel.tcam_mask[1][293][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][294][0]=80'h00000000abf14b53db5d;
sos_loop[0].somModel.tcam_mask[1][294][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][295][0]=80'h00000000d9e701d3b5a1;
sos_loop[0].somModel.tcam_mask[1][295][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][296][0]=80'h00000000ecb4c08dbedf;
sos_loop[0].somModel.tcam_mask[1][296][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][297][0]=80'h0000000059425a4d73e4;
sos_loop[0].somModel.tcam_mask[1][297][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][298][0]=80'h0000000046d500a7b842;
sos_loop[0].somModel.tcam_mask[1][298][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][299][0]=80'h00000000246ba174baea;
sos_loop[0].somModel.tcam_mask[1][299][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][300][0]=80'h00000000e1fa257edda3;
sos_loop[0].somModel.tcam_mask[1][300][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][301][0]=80'h000000009170e9535830;
sos_loop[0].somModel.tcam_mask[1][301][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][302][0]=80'h00000000b0da854090a5;
sos_loop[0].somModel.tcam_mask[1][302][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][303][0]=80'h000000007794a452c0cc;
sos_loop[0].somModel.tcam_mask[1][303][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][304][0]=80'h000000001bb10373944d;
sos_loop[0].somModel.tcam_mask[1][304][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][305][0]=80'h0000000054211c3f4263;
sos_loop[0].somModel.tcam_mask[1][305][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][306][0]=80'h0000000083f85a06a68f;
sos_loop[0].somModel.tcam_mask[1][306][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][307][0]=80'h00000000262df1f69e49;
sos_loop[0].somModel.tcam_mask[1][307][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][308][0]=80'h000000007d107f8ef4a6;
sos_loop[0].somModel.tcam_mask[1][308][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][309][0]=80'h00000000e4475d1bbe07;
sos_loop[0].somModel.tcam_mask[1][309][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][310][0]=80'h00000000f14033c3de26;
sos_loop[0].somModel.tcam_mask[1][310][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][311][0]=80'h000000000eedc1c4b985;
sos_loop[0].somModel.tcam_mask[1][311][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][312][0]=80'h0000000045ea918b6353;
sos_loop[0].somModel.tcam_mask[1][312][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][313][0]=80'h00000000b6e8b1059138;
sos_loop[0].somModel.tcam_mask[1][313][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][314][0]=80'h00000000e2d1f729b709;
sos_loop[0].somModel.tcam_mask[1][314][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][315][0]=80'h000000000358b6eaed36;
sos_loop[0].somModel.tcam_mask[1][315][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[1][316][0]=80'h00000000a67e6c68258f;
sos_loop[0].somModel.tcam_mask[1][316][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][317][0]=80'h000000003aa9c27a9590;
sos_loop[0].somModel.tcam_mask[1][317][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][318][0]=80'h0000000025062337c847;
sos_loop[0].somModel.tcam_mask[1][318][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][319][0]=80'h000000002d9d36fde26f;
sos_loop[0].somModel.tcam_mask[1][319][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][320][0]=80'h00000000a2f4f66c6e72;
sos_loop[0].somModel.tcam_mask[1][320][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][321][0]=80'h00000000d3dbc263b79e;
sos_loop[0].somModel.tcam_mask[1][321][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][322][0]=80'h00000000aa26b833ca5a;
sos_loop[0].somModel.tcam_mask[1][322][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][323][0]=80'h00000000e533d3adc92a;
sos_loop[0].somModel.tcam_mask[1][323][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][324][0]=80'h00000000e7989fff15b9;
sos_loop[0].somModel.tcam_mask[1][324][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][325][0]=80'h00000000204cb109b684;
sos_loop[0].somModel.tcam_mask[1][325][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][326][0]=80'h000000009c86a3258c1c;
sos_loop[0].somModel.tcam_mask[1][326][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][327][0]=80'h0000000033ee6b8cd041;
sos_loop[0].somModel.tcam_mask[1][327][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][328][0]=80'h0000000035cdd2ebe7d4;
sos_loop[0].somModel.tcam_mask[1][328][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][329][0]=80'h00000000fbe9f071ba55;
sos_loop[0].somModel.tcam_mask[1][329][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][330][0]=80'h00000000edbaf396f94d;
sos_loop[0].somModel.tcam_mask[1][330][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][331][0]=80'h000000008f00c6959630;
sos_loop[0].somModel.tcam_mask[1][331][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][332][0]=80'h000000002f0b7d02f677;
sos_loop[0].somModel.tcam_mask[1][332][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][333][0]=80'h0000000084361e779b29;
sos_loop[0].somModel.tcam_mask[1][333][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][334][0]=80'h00000000f9555655c72e;
sos_loop[0].somModel.tcam_mask[1][334][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][335][0]=80'h0000000063fdd2831f64;
sos_loop[0].somModel.tcam_mask[1][335][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][336][0]=80'h0000000044f84811196a;
sos_loop[0].somModel.tcam_mask[1][336][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][337][0]=80'h00000000ee6a7ad1f326;
sos_loop[0].somModel.tcam_mask[1][337][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][338][0]=80'h00000000bd9a0d551dbe;
sos_loop[0].somModel.tcam_mask[1][338][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][339][0]=80'h00000000d77b6743a6d7;
sos_loop[0].somModel.tcam_mask[1][339][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][340][0]=80'h00000000d514be473ad0;
sos_loop[0].somModel.tcam_mask[1][340][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][341][0]=80'h00000000cd8d292c9163;
sos_loop[0].somModel.tcam_mask[1][341][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][342][0]=80'h000000009b96c0a157f3;
sos_loop[0].somModel.tcam_mask[1][342][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][343][0]=80'h000000003990be6ca74b;
sos_loop[0].somModel.tcam_mask[1][343][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][344][0]=80'h00000000878954834a39;
sos_loop[0].somModel.tcam_mask[1][344][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][345][0]=80'h0000000055f55f90aaf2;
sos_loop[0].somModel.tcam_mask[1][345][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][346][0]=80'h000000006528fb359720;
sos_loop[0].somModel.tcam_mask[1][346][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][347][0]=80'h00000000d2e32bd26d81;
sos_loop[0].somModel.tcam_mask[1][347][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][348][0]=80'h000000006cfb0768eaf9;
sos_loop[0].somModel.tcam_mask[1][348][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][349][0]=80'h00000000f605651cbda8;
sos_loop[0].somModel.tcam_mask[1][349][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][350][0]=80'h0000000067afeb283b90;
sos_loop[0].somModel.tcam_mask[1][350][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][351][0]=80'h0000000036956d2c31fd;
sos_loop[0].somModel.tcam_mask[1][351][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][352][0]=80'h00000000eeff5a03dcc4;
sos_loop[0].somModel.tcam_mask[1][352][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][353][0]=80'h0000000068f890ba7165;
sos_loop[0].somModel.tcam_mask[1][353][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][354][0]=80'h00000000859e9ee2a203;
sos_loop[0].somModel.tcam_mask[1][354][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][355][0]=80'h0000000028b1629a2cd1;
sos_loop[0].somModel.tcam_mask[1][355][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][356][0]=80'h00000000f9e13f57f9cb;
sos_loop[0].somModel.tcam_mask[1][356][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][357][0]=80'h000000000eb3232486a6;
sos_loop[0].somModel.tcam_mask[1][357][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][358][0]=80'h00000000812ef34dfa60;
sos_loop[0].somModel.tcam_mask[1][358][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][359][0]=80'h00000000390057c5b93d;
sos_loop[0].somModel.tcam_mask[1][359][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][360][0]=80'h000000009ebf1ea8a8a3;
sos_loop[0].somModel.tcam_mask[1][360][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][361][0]=80'h0000000003511debe665;
sos_loop[0].somModel.tcam_mask[1][361][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[1][362][0]=80'h0000000049fc818617e9;
sos_loop[0].somModel.tcam_mask[1][362][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][363][0]=80'h000000009d37264bcd9f;
sos_loop[0].somModel.tcam_mask[1][363][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][364][0]=80'h000000009a822da69611;
sos_loop[0].somModel.tcam_mask[1][364][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][365][0]=80'h0000000027b44ca01d38;
sos_loop[0].somModel.tcam_mask[1][365][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][366][0]=80'h00000000c0c5608917d4;
sos_loop[0].somModel.tcam_mask[1][366][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][367][0]=80'h0000000081edee6be9a2;
sos_loop[0].somModel.tcam_mask[1][367][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][368][0]=80'h00000000337d2f6ee9f6;
sos_loop[0].somModel.tcam_mask[1][368][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][369][0]=80'h000000003b0f04ce077f;
sos_loop[0].somModel.tcam_mask[1][369][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][370][0]=80'h00000000fde55ff6a820;
sos_loop[0].somModel.tcam_mask[1][370][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][371][0]=80'h00000000dc321bcbeb8f;
sos_loop[0].somModel.tcam_mask[1][371][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][372][0]=80'h000000001bc1c7ca7403;
sos_loop[0].somModel.tcam_mask[1][372][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][373][0]=80'h00000000b7a0d02f7f9a;
sos_loop[0].somModel.tcam_mask[1][373][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][374][0]=80'h000000001c64b4b87959;
sos_loop[0].somModel.tcam_mask[1][374][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][375][0]=80'h000000001e90fcb13925;
sos_loop[0].somModel.tcam_mask[1][375][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][376][0]=80'h000000005ad1dcebe9aa;
sos_loop[0].somModel.tcam_mask[1][376][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][377][0]=80'h0000000045621e9591fb;
sos_loop[0].somModel.tcam_mask[1][377][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][378][0]=80'h0000000059145ef9f8d3;
sos_loop[0].somModel.tcam_mask[1][378][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][379][0]=80'h000000005605b54371f8;
sos_loop[0].somModel.tcam_mask[1][379][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][380][0]=80'h00000000b963e37953dc;
sos_loop[0].somModel.tcam_mask[1][380][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][381][0]=80'h00000000d878910fbeb3;
sos_loop[0].somModel.tcam_mask[1][381][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][382][0]=80'h00000000e8578a861c2c;
sos_loop[0].somModel.tcam_mask[1][382][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][383][0]=80'h000000004ec64f6caae0;
sos_loop[0].somModel.tcam_mask[1][383][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][384][0]=80'h00000000854ba79d2364;
sos_loop[0].somModel.tcam_mask[1][384][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][385][0]=80'h000000002cdf40fd45c7;
sos_loop[0].somModel.tcam_mask[1][385][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][386][0]=80'h00000000a01eaa448072;
sos_loop[0].somModel.tcam_mask[1][386][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][387][0]=80'h00000000d0441435aef0;
sos_loop[0].somModel.tcam_mask[1][387][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][388][0]=80'h000000005d2a8b0aef36;
sos_loop[0].somModel.tcam_mask[1][388][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][389][0]=80'h000000008074ba3f6a36;
sos_loop[0].somModel.tcam_mask[1][389][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][390][0]=80'h000000000053797badc4;
sos_loop[0].somModel.tcam_mask[1][390][0]=80'hffffffffff8000000000;
sos_loop[0].somModel.tcam_data[1][391][0]=80'h000000002ed7fd573cf7;
sos_loop[0].somModel.tcam_mask[1][391][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][392][0]=80'h00000000e5883e982b3c;
sos_loop[0].somModel.tcam_mask[1][392][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][393][0]=80'h0000000053a2748e29f6;
sos_loop[0].somModel.tcam_mask[1][393][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][394][0]=80'h000000005ca1a2544aa9;
sos_loop[0].somModel.tcam_mask[1][394][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][395][0]=80'h00000000e3f9ded7caed;
sos_loop[0].somModel.tcam_mask[1][395][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][396][0]=80'h00000000a3643184f60a;
sos_loop[0].somModel.tcam_mask[1][396][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][397][0]=80'h000000002852f1edb5fa;
sos_loop[0].somModel.tcam_mask[1][397][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][398][0]=80'h000000003244642a522c;
sos_loop[0].somModel.tcam_mask[1][398][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][399][0]=80'h00000000577ae1143ac3;
sos_loop[0].somModel.tcam_mask[1][399][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][400][0]=80'h00000000d116b38ae558;
sos_loop[0].somModel.tcam_mask[1][400][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][401][0]=80'h00000000ef6f5c21938c;
sos_loop[0].somModel.tcam_mask[1][401][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][402][0]=80'h00000000c7ae9723534c;
sos_loop[0].somModel.tcam_mask[1][402][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][403][0]=80'h0000000012ee7fec5c3e;
sos_loop[0].somModel.tcam_mask[1][403][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][404][0]=80'h000000008ceb8fe138f0;
sos_loop[0].somModel.tcam_mask[1][404][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][405][0]=80'h00000000ac6c00b6a8d2;
sos_loop[0].somModel.tcam_mask[1][405][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][406][0]=80'h00000000b15acb7a407c;
sos_loop[0].somModel.tcam_mask[1][406][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][407][0]=80'h00000000fe01162b7c3d;
sos_loop[0].somModel.tcam_mask[1][407][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][408][0]=80'h000000003ca520daccf9;
sos_loop[0].somModel.tcam_mask[1][408][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][409][0]=80'h000000001ddba06c2730;
sos_loop[0].somModel.tcam_mask[1][409][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][410][0]=80'h000000008c25018e78c8;
sos_loop[0].somModel.tcam_mask[1][410][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][411][0]=80'h00000000294e58af58b8;
sos_loop[0].somModel.tcam_mask[1][411][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][412][0]=80'h0000000025431f6f1ca8;
sos_loop[0].somModel.tcam_mask[1][412][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][413][0]=80'h000000000d4e0d35b1bb;
sos_loop[0].somModel.tcam_mask[1][413][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][414][0]=80'h00000000288f8de89002;
sos_loop[0].somModel.tcam_mask[1][414][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][415][0]=80'h00000000bbd2142468fd;
sos_loop[0].somModel.tcam_mask[1][415][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][416][0]=80'h000000009285b15180ce;
sos_loop[0].somModel.tcam_mask[1][416][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][417][0]=80'h0000000089d7c1092a1f;
sos_loop[0].somModel.tcam_mask[1][417][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][418][0]=80'h00000000bc5113c19cfc;
sos_loop[0].somModel.tcam_mask[1][418][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][419][0]=80'h00000000cb0ad767c3ff;
sos_loop[0].somModel.tcam_mask[1][419][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][420][0]=80'h0000000064d3dedd3b11;
sos_loop[0].somModel.tcam_mask[1][420][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][421][0]=80'h000000001e5eb38233fd;
sos_loop[0].somModel.tcam_mask[1][421][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][422][0]=80'h00000000d9b98809ae51;
sos_loop[0].somModel.tcam_mask[1][422][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][423][0]=80'h000000005f3093fd17e5;
sos_loop[0].somModel.tcam_mask[1][423][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][424][0]=80'h000000008f220f87bb88;
sos_loop[0].somModel.tcam_mask[1][424][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][425][0]=80'h000000002effec1166ca;
sos_loop[0].somModel.tcam_mask[1][425][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][426][0]=80'h000000008efae6f79380;
sos_loop[0].somModel.tcam_mask[1][426][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][427][0]=80'h000000001e1735b714f1;
sos_loop[0].somModel.tcam_mask[1][427][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][428][0]=80'h0000000074b95b6a5e36;
sos_loop[0].somModel.tcam_mask[1][428][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][429][0]=80'h00000000ad17df6d5280;
sos_loop[0].somModel.tcam_mask[1][429][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][430][0]=80'h00000000d9cc5ca6a92a;
sos_loop[0].somModel.tcam_mask[1][430][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][431][0]=80'h00000000bcc4cdb632c7;
sos_loop[0].somModel.tcam_mask[1][431][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][432][0]=80'h0000000078702dc7b992;
sos_loop[0].somModel.tcam_mask[1][432][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][433][0]=80'h000000004c0ae5cc4065;
sos_loop[0].somModel.tcam_mask[1][433][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][434][0]=80'h000000006d192447580c;
sos_loop[0].somModel.tcam_mask[1][434][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][435][0]=80'h000000004082eb1df830;
sos_loop[0].somModel.tcam_mask[1][435][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][436][0]=80'h000000006789fbb57be3;
sos_loop[0].somModel.tcam_mask[1][436][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][437][0]=80'h00000000271e20654263;
sos_loop[0].somModel.tcam_mask[1][437][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][438][0]=80'h0000000046c0f48c2876;
sos_loop[0].somModel.tcam_mask[1][438][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][439][0]=80'h00000000b0e588475012;
sos_loop[0].somModel.tcam_mask[1][439][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][440][0]=80'h00000000f3bd582ea928;
sos_loop[0].somModel.tcam_mask[1][440][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][441][0]=80'h000000002138e3a06726;
sos_loop[0].somModel.tcam_mask[1][441][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][442][0]=80'h00000000a916c7e72f2c;
sos_loop[0].somModel.tcam_mask[1][442][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][443][0]=80'h00000000b731cb59fe72;
sos_loop[0].somModel.tcam_mask[1][443][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][444][0]=80'h00000000abcdc1e96b29;
sos_loop[0].somModel.tcam_mask[1][444][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][445][0]=80'h0000000038bcc2b05d26;
sos_loop[0].somModel.tcam_mask[1][445][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][446][0]=80'h0000000013f98cd1dbbd;
sos_loop[0].somModel.tcam_mask[1][446][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][447][0]=80'h00000000e592927a0a89;
sos_loop[0].somModel.tcam_mask[1][447][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][448][0]=80'h000000009470cfe0bd38;
sos_loop[0].somModel.tcam_mask[1][448][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][449][0]=80'h00000000ab62ba7b123c;
sos_loop[0].somModel.tcam_mask[1][449][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][450][0]=80'h00000000c9793372f335;
sos_loop[0].somModel.tcam_mask[1][450][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][451][0]=80'h0000000017c05008dfd2;
sos_loop[0].somModel.tcam_mask[1][451][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][452][0]=80'h000000007938cdcbad6d;
sos_loop[0].somModel.tcam_mask[1][452][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][453][0]=80'h00000000282455e8a649;
sos_loop[0].somModel.tcam_mask[1][453][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][454][0]=80'h00000000d4b10f962ebd;
sos_loop[0].somModel.tcam_mask[1][454][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][455][0]=80'h00000000ee2a158883b5;
sos_loop[0].somModel.tcam_mask[1][455][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][456][0]=80'h00000000906a9ad30087;
sos_loop[0].somModel.tcam_mask[1][456][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][457][0]=80'h0000000004282827d137;
sos_loop[0].somModel.tcam_mask[1][457][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[1][458][0]=80'h00000000585a643eec07;
sos_loop[0].somModel.tcam_mask[1][458][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][459][0]=80'h00000000eb073e9ed5c7;
sos_loop[0].somModel.tcam_mask[1][459][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][460][0]=80'h00000000021b4376f56e;
sos_loop[0].somModel.tcam_mask[1][460][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[1][461][0]=80'h00000000bd2b7e328666;
sos_loop[0].somModel.tcam_mask[1][461][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][462][0]=80'h00000000f6b6101e438d;
sos_loop[0].somModel.tcam_mask[1][462][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][463][0]=80'h00000000908022cd936f;
sos_loop[0].somModel.tcam_mask[1][463][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][464][0]=80'h000000007511ee9fa2de;
sos_loop[0].somModel.tcam_mask[1][464][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][465][0]=80'h00000000374776fb63b1;
sos_loop[0].somModel.tcam_mask[1][465][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][466][0]=80'h00000000d65c8503efa5;
sos_loop[0].somModel.tcam_mask[1][466][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][467][0]=80'h000000009ad572e1b926;
sos_loop[0].somModel.tcam_mask[1][467][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][468][0]=80'h000000009e796c3e4446;
sos_loop[0].somModel.tcam_mask[1][468][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][469][0]=80'h0000000081296115c65e;
sos_loop[0].somModel.tcam_mask[1][469][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][470][0]=80'h000000002ef37672dd00;
sos_loop[0].somModel.tcam_mask[1][470][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][471][0]=80'h000000001be09a9632b7;
sos_loop[0].somModel.tcam_mask[1][471][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][472][0]=80'h00000000a0251ac3bdd7;
sos_loop[0].somModel.tcam_mask[1][472][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][473][0]=80'h00000000fa7f865e62ee;
sos_loop[0].somModel.tcam_mask[1][473][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][474][0]=80'h00000000290b9b7a1e05;
sos_loop[0].somModel.tcam_mask[1][474][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][475][0]=80'h000000007f8e37e50737;
sos_loop[0].somModel.tcam_mask[1][475][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][476][0]=80'h00000000e96a1056fbe0;
sos_loop[0].somModel.tcam_mask[1][476][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][477][0]=80'h00000000492b7df8136d;
sos_loop[0].somModel.tcam_mask[1][477][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][478][0]=80'h00000000b391bb6cff61;
sos_loop[0].somModel.tcam_mask[1][478][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][479][0]=80'h00000000b82153980608;
sos_loop[0].somModel.tcam_mask[1][479][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][480][0]=80'h00000000abcbdbe195e1;
sos_loop[0].somModel.tcam_mask[1][480][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][481][0]=80'h00000000fcefb0d3fb08;
sos_loop[0].somModel.tcam_mask[1][481][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][482][0]=80'h00000000789711b0a797;
sos_loop[0].somModel.tcam_mask[1][482][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][483][0]=80'h000000005cf2068e30a7;
sos_loop[0].somModel.tcam_mask[1][483][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][484][0]=80'h00000000d4dfd545d947;
sos_loop[0].somModel.tcam_mask[1][484][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][485][0]=80'h000000004926b200a921;
sos_loop[0].somModel.tcam_mask[1][485][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][486][0]=80'h00000000c373a403d24b;
sos_loop[0].somModel.tcam_mask[1][486][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][487][0]=80'h000000007e109be15c54;
sos_loop[0].somModel.tcam_mask[1][487][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][488][0]=80'h00000000b79c76af4364;
sos_loop[0].somModel.tcam_mask[1][488][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][489][0]=80'h0000000042ad91b91308;
sos_loop[0].somModel.tcam_mask[1][489][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][490][0]=80'h00000000923c87528181;
sos_loop[0].somModel.tcam_mask[1][490][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][491][0]=80'h000000006927aecffc09;
sos_loop[0].somModel.tcam_mask[1][491][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][492][0]=80'h00000000b0d09ccc302d;
sos_loop[0].somModel.tcam_mask[1][492][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][493][0]=80'h00000000a4234997ebd8;
sos_loop[0].somModel.tcam_mask[1][493][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][494][0]=80'h000000001ed04fa1ec97;
sos_loop[0].somModel.tcam_mask[1][494][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][495][0]=80'h000000009892ee4621b6;
sos_loop[0].somModel.tcam_mask[1][495][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][496][0]=80'h00000000cfc813360aaa;
sos_loop[0].somModel.tcam_mask[1][496][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][497][0]=80'h000000005e383a86df15;
sos_loop[0].somModel.tcam_mask[1][497][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][498][0]=80'h00000000975c188f1dbe;
sos_loop[0].somModel.tcam_mask[1][498][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][499][0]=80'h000000005ae15f494a6f;
sos_loop[0].somModel.tcam_mask[1][499][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][500][0]=80'h00000000ba60c9b84434;
sos_loop[0].somModel.tcam_mask[1][500][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][501][0]=80'h00000000ec5378e383d8;
sos_loop[0].somModel.tcam_mask[1][501][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][502][0]=80'h00000000c6f584a0c437;
sos_loop[0].somModel.tcam_mask[1][502][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][503][0]=80'h0000000037b198167e84;
sos_loop[0].somModel.tcam_mask[1][503][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][504][0]=80'h00000000d5a720e74827;
sos_loop[0].somModel.tcam_mask[1][504][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][505][0]=80'h0000000002b27ae1774a;
sos_loop[0].somModel.tcam_mask[1][505][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[1][506][0]=80'h00000000d7ccbf2c8a33;
sos_loop[0].somModel.tcam_mask[1][506][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][507][0]=80'h00000000d7821106381a;
sos_loop[0].somModel.tcam_mask[1][507][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][508][0]=80'h0000000027abf231a4f3;
sos_loop[0].somModel.tcam_mask[1][508][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][509][0]=80'h00000000f6b0f88997b0;
sos_loop[0].somModel.tcam_mask[1][509][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][510][0]=80'h000000008bf13cd9575c;
sos_loop[0].somModel.tcam_mask[1][510][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][511][0]=80'h000000003269043ae182;
sos_loop[0].somModel.tcam_mask[1][511][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][512][0]=80'h00000000a08b34cab3ff;
sos_loop[0].somModel.tcam_mask[1][512][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][513][0]=80'h0000000035f72570ae87;
sos_loop[0].somModel.tcam_mask[1][513][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][514][0]=80'h00000000ef37fd8baffb;
sos_loop[0].somModel.tcam_mask[1][514][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][515][0]=80'h00000000caff585f4b5f;
sos_loop[0].somModel.tcam_mask[1][515][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][516][0]=80'h0000000076eee9f3d2c5;
sos_loop[0].somModel.tcam_mask[1][516][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][517][0]=80'h00000000af06beec59cb;
sos_loop[0].somModel.tcam_mask[1][517][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][518][0]=80'h0000000082c90775e233;
sos_loop[0].somModel.tcam_mask[1][518][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][519][0]=80'h00000000fe0847448447;
sos_loop[0].somModel.tcam_mask[1][519][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][520][0]=80'h00000000f0cb1f28c22a;
sos_loop[0].somModel.tcam_mask[1][520][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][521][0]=80'h000000007079f2078cc4;
sos_loop[0].somModel.tcam_mask[1][521][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][522][0]=80'h000000006abd25be785f;
sos_loop[0].somModel.tcam_mask[1][522][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][523][0]=80'h00000000dfdfc2f15c4d;
sos_loop[0].somModel.tcam_mask[1][523][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][524][0]=80'h00000000c9d15a930997;
sos_loop[0].somModel.tcam_mask[1][524][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][525][0]=80'h00000000a894e1e563f1;
sos_loop[0].somModel.tcam_mask[1][525][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][526][0]=80'h00000000a964fe119d5f;
sos_loop[0].somModel.tcam_mask[1][526][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][527][0]=80'h000000009dafde935b53;
sos_loop[0].somModel.tcam_mask[1][527][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][528][0]=80'h000000000e906f4b5764;
sos_loop[0].somModel.tcam_mask[1][528][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][529][0]=80'h00000000216048dbe8e2;
sos_loop[0].somModel.tcam_mask[1][529][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][530][0]=80'h00000000c08f3732c7eb;
sos_loop[0].somModel.tcam_mask[1][530][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][531][0]=80'h00000000b72142bca4aa;
sos_loop[0].somModel.tcam_mask[1][531][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][532][0]=80'h0000000067a2ce8a5e0e;
sos_loop[0].somModel.tcam_mask[1][532][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][533][0]=80'h000000005819e54162b8;
sos_loop[0].somModel.tcam_mask[1][533][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][534][0]=80'h00000000f81fb7436abb;
sos_loop[0].somModel.tcam_mask[1][534][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][535][0]=80'h0000000031d8f5200247;
sos_loop[0].somModel.tcam_mask[1][535][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][536][0]=80'h00000000607df517446f;
sos_loop[0].somModel.tcam_mask[1][536][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][537][0]=80'h000000009501b95b8eee;
sos_loop[0].somModel.tcam_mask[1][537][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][538][0]=80'h000000004ac80e1571f3;
sos_loop[0].somModel.tcam_mask[1][538][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][539][0]=80'h00000000397eabef6f73;
sos_loop[0].somModel.tcam_mask[1][539][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][540][0]=80'h0000000058330b72f740;
sos_loop[0].somModel.tcam_mask[1][540][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][541][0]=80'h00000000b091099c5208;
sos_loop[0].somModel.tcam_mask[1][541][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][542][0]=80'h000000008c922af3d544;
sos_loop[0].somModel.tcam_mask[1][542][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][543][0]=80'h000000001ef54a94a1aa;
sos_loop[0].somModel.tcam_mask[1][543][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][544][0]=80'h00000000eafb610d3307;
sos_loop[0].somModel.tcam_mask[1][544][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][545][0]=80'h000000008f6e4315ccf3;
sos_loop[0].somModel.tcam_mask[1][545][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][546][0]=80'h00000000be335ca6def9;
sos_loop[0].somModel.tcam_mask[1][546][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][547][0]=80'h00000000ee0d6e2944d0;
sos_loop[0].somModel.tcam_mask[1][547][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][548][0]=80'h000000000f79f7b4fbc4;
sos_loop[0].somModel.tcam_mask[1][548][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][549][0]=80'h0000000016a4b9b11745;
sos_loop[0].somModel.tcam_mask[1][549][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][550][0]=80'h00000000b854815e349a;
sos_loop[0].somModel.tcam_mask[1][550][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][551][0]=80'h000000008264f4b38d53;
sos_loop[0].somModel.tcam_mask[1][551][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][552][0]=80'h0000000002b31497dfe4;
sos_loop[0].somModel.tcam_mask[1][552][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[1][553][0]=80'h000000003874850e3664;
sos_loop[0].somModel.tcam_mask[1][553][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][554][0]=80'h000000001e03504fc71e;
sos_loop[0].somModel.tcam_mask[1][554][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][555][0]=80'h00000000ac17c1eed961;
sos_loop[0].somModel.tcam_mask[1][555][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][556][0]=80'h000000008b4a08190ea6;
sos_loop[0].somModel.tcam_mask[1][556][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][557][0]=80'h000000001a089420fe6b;
sos_loop[0].somModel.tcam_mask[1][557][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][558][0]=80'h00000000db0519d32d54;
sos_loop[0].somModel.tcam_mask[1][558][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][559][0]=80'h00000000d606b6890ccf;
sos_loop[0].somModel.tcam_mask[1][559][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][560][0]=80'h000000003a30d200a52e;
sos_loop[0].somModel.tcam_mask[1][560][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][561][0]=80'h00000000e1d629596d55;
sos_loop[0].somModel.tcam_mask[1][561][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][562][0]=80'h0000000059f8bd5018fa;
sos_loop[0].somModel.tcam_mask[1][562][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][563][0]=80'h0000000018c7b4420188;
sos_loop[0].somModel.tcam_mask[1][563][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][564][0]=80'h00000000381e1bed184a;
sos_loop[0].somModel.tcam_mask[1][564][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][565][0]=80'h00000000d4a5ae2c135b;
sos_loop[0].somModel.tcam_mask[1][565][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][566][0]=80'h00000000e97961ccdcd0;
sos_loop[0].somModel.tcam_mask[1][566][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][567][0]=80'h00000000737a13e21630;
sos_loop[0].somModel.tcam_mask[1][567][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][568][0]=80'h000000006576d31493a8;
sos_loop[0].somModel.tcam_mask[1][568][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][569][0]=80'h0000000016d47d0405e3;
sos_loop[0].somModel.tcam_mask[1][569][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][570][0]=80'h0000000033d13d02eaa0;
sos_loop[0].somModel.tcam_mask[1][570][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][571][0]=80'h00000000d7950dbecaa4;
sos_loop[0].somModel.tcam_mask[1][571][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][572][0]=80'h0000000058f7de01221a;
sos_loop[0].somModel.tcam_mask[1][572][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][573][0]=80'h00000000f297721ec69a;
sos_loop[0].somModel.tcam_mask[1][573][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][574][0]=80'h00000000fa8073a2c40f;
sos_loop[0].somModel.tcam_mask[1][574][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][575][0]=80'h00000000991dda905a7c;
sos_loop[0].somModel.tcam_mask[1][575][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][576][0]=80'h00000000b81a5d03ce28;
sos_loop[0].somModel.tcam_mask[1][576][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][577][0]=80'h00000000793b9c78b761;
sos_loop[0].somModel.tcam_mask[1][577][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][578][0]=80'h00000000048d383e9db0;
sos_loop[0].somModel.tcam_mask[1][578][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[1][579][0]=80'h0000000094a5e12a8d29;
sos_loop[0].somModel.tcam_mask[1][579][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][580][0]=80'h0000000057351e593cda;
sos_loop[0].somModel.tcam_mask[1][580][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][581][0]=80'h0000000087cf3b2441aa;
sos_loop[0].somModel.tcam_mask[1][581][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][582][0]=80'h00000000f43a10956f47;
sos_loop[0].somModel.tcam_mask[1][582][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][583][0]=80'h00000000de3fb55a35c3;
sos_loop[0].somModel.tcam_mask[1][583][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][584][0]=80'h000000008018c8ac27bd;
sos_loop[0].somModel.tcam_mask[1][584][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][585][0]=80'h000000005a5c46dda87a;
sos_loop[0].somModel.tcam_mask[1][585][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][586][0]=80'h000000003c0309aa8715;
sos_loop[0].somModel.tcam_mask[1][586][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][587][0]=80'h0000000068918363bb53;
sos_loop[0].somModel.tcam_mask[1][587][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][588][0]=80'h000000001a50f7d56556;
sos_loop[0].somModel.tcam_mask[1][588][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][589][0]=80'h000000004141bcc97dea;
sos_loop[0].somModel.tcam_mask[1][589][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][590][0]=80'h0000000030b786d0937c;
sos_loop[0].somModel.tcam_mask[1][590][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][591][0]=80'h000000004a0defcfa63e;
sos_loop[0].somModel.tcam_mask[1][591][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][592][0]=80'h000000004fefa8a8325b;
sos_loop[0].somModel.tcam_mask[1][592][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][593][0]=80'h0000000065be949c2999;
sos_loop[0].somModel.tcam_mask[1][593][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][594][0]=80'h00000000e228f54db17f;
sos_loop[0].somModel.tcam_mask[1][594][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][595][0]=80'h00000000ded2a0f4626e;
sos_loop[0].somModel.tcam_mask[1][595][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][596][0]=80'h0000000043be668ec635;
sos_loop[0].somModel.tcam_mask[1][596][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][597][0]=80'h00000000642c6fad96e2;
sos_loop[0].somModel.tcam_mask[1][597][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][598][0]=80'h00000000869bf468988e;
sos_loop[0].somModel.tcam_mask[1][598][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][599][0]=80'h00000000423d784e463c;
sos_loop[0].somModel.tcam_mask[1][599][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][600][0]=80'h000000009e0d7122e5d0;
sos_loop[0].somModel.tcam_mask[1][600][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][601][0]=80'h000000000bbf5f3f9a3d;
sos_loop[0].somModel.tcam_mask[1][601][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][602][0]=80'h000000004d41bb7e83d4;
sos_loop[0].somModel.tcam_mask[1][602][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][603][0]=80'h0000000009fe21480bf2;
sos_loop[0].somModel.tcam_mask[1][603][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][604][0]=80'h000000002daa4544c73c;
sos_loop[0].somModel.tcam_mask[1][604][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][605][0]=80'h00000000de9abc1ba70d;
sos_loop[0].somModel.tcam_mask[1][605][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][606][0]=80'h0000000074b4b8faa3cd;
sos_loop[0].somModel.tcam_mask[1][606][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][607][0]=80'h0000000053ffaa95bde0;
sos_loop[0].somModel.tcam_mask[1][607][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][608][0]=80'h000000007626b2b6c686;
sos_loop[0].somModel.tcam_mask[1][608][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][609][0]=80'h0000000063c350b895ee;
sos_loop[0].somModel.tcam_mask[1][609][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][610][0]=80'h00000000f4023a42fb3d;
sos_loop[0].somModel.tcam_mask[1][610][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][611][0]=80'h00000000d063b376df50;
sos_loop[0].somModel.tcam_mask[1][611][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][612][0]=80'h00000000ef9c58730d40;
sos_loop[0].somModel.tcam_mask[1][612][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][613][0]=80'h00000000b7f07d70beeb;
sos_loop[0].somModel.tcam_mask[1][613][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][614][0]=80'h00000000c6e6e5c33fca;
sos_loop[0].somModel.tcam_mask[1][614][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][615][0]=80'h0000000032388657a2c4;
sos_loop[0].somModel.tcam_mask[1][615][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][616][0]=80'h000000006714ee2ee494;
sos_loop[0].somModel.tcam_mask[1][616][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][617][0]=80'h0000000095e542ea9383;
sos_loop[0].somModel.tcam_mask[1][617][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][618][0]=80'h000000006ee62d6a2974;
sos_loop[0].somModel.tcam_mask[1][618][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][619][0]=80'h00000000992d98d8c860;
sos_loop[0].somModel.tcam_mask[1][619][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][620][0]=80'h000000009d01df2dd16f;
sos_loop[0].somModel.tcam_mask[1][620][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][621][0]=80'h00000000529561ddc2c7;
sos_loop[0].somModel.tcam_mask[1][621][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][622][0]=80'h00000000ed170481df56;
sos_loop[0].somModel.tcam_mask[1][622][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][623][0]=80'h000000008053bfce2d39;
sos_loop[0].somModel.tcam_mask[1][623][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][624][0]=80'h000000002b3565e41eba;
sos_loop[0].somModel.tcam_mask[1][624][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][625][0]=80'h00000000d039014a8676;
sos_loop[0].somModel.tcam_mask[1][625][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][626][0]=80'h000000008aead6f8e415;
sos_loop[0].somModel.tcam_mask[1][626][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][627][0]=80'h00000000bc559f92bfc8;
sos_loop[0].somModel.tcam_mask[1][627][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][628][0]=80'h000000009ef7759a4335;
sos_loop[0].somModel.tcam_mask[1][628][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][629][0]=80'h0000000036050c4a38da;
sos_loop[0].somModel.tcam_mask[1][629][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][630][0]=80'h000000003a029f298309;
sos_loop[0].somModel.tcam_mask[1][630][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][631][0]=80'h00000000c13120cb0493;
sos_loop[0].somModel.tcam_mask[1][631][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][632][0]=80'h000000004a807d566fcc;
sos_loop[0].somModel.tcam_mask[1][632][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][633][0]=80'h00000000f4264c62ed60;
sos_loop[0].somModel.tcam_mask[1][633][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][634][0]=80'h0000000060c439a2621c;
sos_loop[0].somModel.tcam_mask[1][634][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][635][0]=80'h0000000066b493e0fe24;
sos_loop[0].somModel.tcam_mask[1][635][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][636][0]=80'h000000009b6927b93f7d;
sos_loop[0].somModel.tcam_mask[1][636][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][637][0]=80'h00000000704b7af77695;
sos_loop[0].somModel.tcam_mask[1][637][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][638][0]=80'h0000000040ab28bca25f;
sos_loop[0].somModel.tcam_mask[1][638][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][639][0]=80'h00000000c17bb0702ae1;
sos_loop[0].somModel.tcam_mask[1][639][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][640][0]=80'h00000000b0d05cb346d2;
sos_loop[0].somModel.tcam_mask[1][640][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][641][0]=80'h00000000cb0be3f40df1;
sos_loop[0].somModel.tcam_mask[1][641][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][642][0]=80'h00000000b40e6c1f67e0;
sos_loop[0].somModel.tcam_mask[1][642][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][643][0]=80'h00000000dd08373eb7e2;
sos_loop[0].somModel.tcam_mask[1][643][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][644][0]=80'h00000000321f38e6c645;
sos_loop[0].somModel.tcam_mask[1][644][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][645][0]=80'h00000000022f54ffa712;
sos_loop[0].somModel.tcam_mask[1][645][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[1][646][0]=80'h00000000175711491a12;
sos_loop[0].somModel.tcam_mask[1][646][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][647][0]=80'h000000005c4334e83dbf;
sos_loop[0].somModel.tcam_mask[1][647][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][648][0]=80'h000000007401586b796c;
sos_loop[0].somModel.tcam_mask[1][648][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][649][0]=80'h000000001064da257814;
sos_loop[0].somModel.tcam_mask[1][649][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][650][0]=80'h0000000033aa97849759;
sos_loop[0].somModel.tcam_mask[1][650][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][651][0]=80'h00000000dd749f6d10f2;
sos_loop[0].somModel.tcam_mask[1][651][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][652][0]=80'h0000000032ec91b393dd;
sos_loop[0].somModel.tcam_mask[1][652][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][653][0]=80'h0000000014cc9cebd56f;
sos_loop[0].somModel.tcam_mask[1][653][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][654][0]=80'h00000000fa1a640d3120;
sos_loop[0].somModel.tcam_mask[1][654][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][655][0]=80'h00000000f4e3f6a941f0;
sos_loop[0].somModel.tcam_mask[1][655][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][656][0]=80'h00000000d00f18748035;
sos_loop[0].somModel.tcam_mask[1][656][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][657][0]=80'h00000000471f97f6e335;
sos_loop[0].somModel.tcam_mask[1][657][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][658][0]=80'h0000000025d72449c9e0;
sos_loop[0].somModel.tcam_mask[1][658][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][659][0]=80'h0000000054f6d49980a3;
sos_loop[0].somModel.tcam_mask[1][659][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][660][0]=80'h00000000d9a3a9015e31;
sos_loop[0].somModel.tcam_mask[1][660][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][661][0]=80'h000000007ca54a31df80;
sos_loop[0].somModel.tcam_mask[1][661][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][662][0]=80'h000000002727fd6cbcb5;
sos_loop[0].somModel.tcam_mask[1][662][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][663][0]=80'h000000008d849e8d0bd6;
sos_loop[0].somModel.tcam_mask[1][663][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][664][0]=80'h00000000c7917e2857fc;
sos_loop[0].somModel.tcam_mask[1][664][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][665][0]=80'h00000000c114d4bda130;
sos_loop[0].somModel.tcam_mask[1][665][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][666][0]=80'h000000000be6a2e10c1a;
sos_loop[0].somModel.tcam_mask[1][666][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][667][0]=80'h00000000ef3b11cfca80;
sos_loop[0].somModel.tcam_mask[1][667][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][668][0]=80'h00000000da6802e720b7;
sos_loop[0].somModel.tcam_mask[1][668][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][669][0]=80'h00000000b955999acc64;
sos_loop[0].somModel.tcam_mask[1][669][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][670][0]=80'h000000000dc76ebecea5;
sos_loop[0].somModel.tcam_mask[1][670][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][671][0]=80'h000000003d59e483ea45;
sos_loop[0].somModel.tcam_mask[1][671][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][672][0]=80'h000000008e98064d1c2c;
sos_loop[0].somModel.tcam_mask[1][672][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][673][0]=80'h00000000111c13b657b7;
sos_loop[0].somModel.tcam_mask[1][673][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[1][674][0]=80'h00000000ef7d1553096c;
sos_loop[0].somModel.tcam_mask[1][674][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][675][0]=80'h0000000091047a599dcf;
sos_loop[0].somModel.tcam_mask[1][675][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][676][0]=80'h00000000a8423d3eddb2;
sos_loop[0].somModel.tcam_mask[1][676][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][677][0]=80'h000000000cfd34e86e5f;
sos_loop[0].somModel.tcam_mask[1][677][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[1][678][0]=80'h0000000075ebdb494049;
sos_loop[0].somModel.tcam_mask[1][678][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][679][0]=80'h000000003b3640c4d206;
sos_loop[0].somModel.tcam_mask[1][679][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][680][0]=80'h00000000d119b635c7bc;
sos_loop[0].somModel.tcam_mask[1][680][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][681][0]=80'h00000000719073427062;
sos_loop[0].somModel.tcam_mask[1][681][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][682][0]=80'h000000005d2633c1c0c6;
sos_loop[0].somModel.tcam_mask[1][682][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][683][0]=80'h000000005ffe5556f980;
sos_loop[0].somModel.tcam_mask[1][683][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][684][0]=80'h0000000061e8d059e1f9;
sos_loop[0].somModel.tcam_mask[1][684][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][685][0]=80'h00000000203ef10ced3e;
sos_loop[0].somModel.tcam_mask[1][685][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][686][0]=80'h000000009eee630d6efc;
sos_loop[0].somModel.tcam_mask[1][686][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][687][0]=80'h000000006322298a3a7b;
sos_loop[0].somModel.tcam_mask[1][687][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][688][0]=80'h00000000f40c4bfc22fa;
sos_loop[0].somModel.tcam_mask[1][688][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][689][0]=80'h00000000fa5c7b97f665;
sos_loop[0].somModel.tcam_mask[1][689][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][690][0]=80'h00000000ef9dfeb948eb;
sos_loop[0].somModel.tcam_mask[1][690][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][691][0]=80'h00000000382de4729315;
sos_loop[0].somModel.tcam_mask[1][691][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][692][0]=80'h0000000045bb0fa48950;
sos_loop[0].somModel.tcam_mask[1][692][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][693][0]=80'h000000002ab5c380b341;
sos_loop[0].somModel.tcam_mask[1][693][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[1][694][0]=80'h000000009f6273d1e971;
sos_loop[0].somModel.tcam_mask[1][694][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][695][0]=80'h00000000bc88ff2fe271;
sos_loop[0].somModel.tcam_mask[1][695][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][696][0]=80'h00000000c345fbecc076;
sos_loop[0].somModel.tcam_mask[1][696][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][697][0]=80'h00000000b6b2b6a8914d;
sos_loop[0].somModel.tcam_mask[1][697][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][698][0]=80'h0000000069611d6f9e84;
sos_loop[0].somModel.tcam_mask[1][698][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[1][699][0]=80'h00000000bb21e0ea60b7;
sos_loop[0].somModel.tcam_mask[1][699][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[1][700][0]=80'h00000000247897856c97;
sos_loop[0].somModel.tcam_mask[1][700][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.sram_dat[1][0][0]=96'hdeadbf;
sos_loop[0].somModel.sram_ptr[1][0]=939;
sos_loop[0].somModel.sram_dat[1][1][0]=96'h93d46a;
sos_loop[0].somModel.sram_ptr[1][1]=2;
sos_loop[0].somModel.sram_dat[1][2][0]=96'hd2356f;
sos_loop[0].somModel.sram_ptr[1][2]=2;
sos_loop[0].somModel.sram_dat[1][3][0]=96'h676259;
sos_loop[0].somModel.sram_ptr[1][3]=2;
sos_loop[0].somModel.sram_dat[1][4][0]=96'h46079b;
sos_loop[0].somModel.sram_ptr[1][4]=2;
sos_loop[0].somModel.sram_dat[1][5][0]=96'h8c8892;
sos_loop[0].somModel.sram_ptr[1][5]=2;
sos_loop[0].somModel.sram_dat[1][6][0]=96'h17cf44;
sos_loop[0].somModel.sram_ptr[1][6]=2;
sos_loop[0].somModel.sram_dat[1][7][0]=96'hbc724b;
sos_loop[0].somModel.sram_ptr[1][7]=2;
sos_loop[0].somModel.sram_dat[1][8][0]=96'he97981;
sos_loop[0].somModel.sram_ptr[1][8]=2;
sos_loop[0].somModel.sram_dat[1][9][0]=96'h77a9de;
sos_loop[0].somModel.sram_ptr[1][9]=2;
sos_loop[0].somModel.sram_dat[1][10][0]=96'h2b7a6c;
sos_loop[0].somModel.sram_ptr[1][10]=2;
sos_loop[0].somModel.sram_dat[1][11][0]=96'h504864;
sos_loop[0].somModel.sram_ptr[1][11]=2;
sos_loop[0].somModel.sram_dat[1][12][0]=96'h8c6bb5;
sos_loop[0].somModel.sram_ptr[1][12]=2;
sos_loop[0].somModel.sram_dat[1][13][0]=96'h7afada;
sos_loop[0].somModel.sram_ptr[1][13]=2;
sos_loop[0].somModel.sram_dat[1][14][0]=96'hcc3650;
sos_loop[0].somModel.sram_ptr[1][14]=2;
sos_loop[0].somModel.sram_dat[1][15][0]=96'hdde1;
sos_loop[0].somModel.sram_ptr[1][15]=2;
sos_loop[0].somModel.sram_dat[1][16][0]=96'h41bae2;
sos_loop[0].somModel.sram_ptr[1][16]=2;
sos_loop[0].somModel.sram_dat[1][17][0]=96'h4b4f80;
sos_loop[0].somModel.sram_ptr[1][17]=2;
sos_loop[0].somModel.sram_dat[1][18][0]=96'hccad23;
sos_loop[0].somModel.sram_ptr[1][18]=2;
sos_loop[0].somModel.sram_dat[1][19][0]=96'h987d18;
sos_loop[0].somModel.sram_ptr[1][19]=2;
sos_loop[0].somModel.sram_dat[1][20][0]=96'h354214;
sos_loop[0].somModel.sram_ptr[1][20]=2;
sos_loop[0].somModel.sram_dat[1][21][0]=96'h1b5bf0;
sos_loop[0].somModel.sram_ptr[1][21]=2;
sos_loop[0].somModel.sram_dat[1][22][0]=96'hcfcfe0;
sos_loop[0].somModel.sram_ptr[1][22]=2;
sos_loop[0].somModel.sram_dat[1][23][0]=96'h5dfdd7;
sos_loop[0].somModel.sram_ptr[1][23]=2;
sos_loop[0].somModel.sram_dat[1][24][0]=96'hf65193;
sos_loop[0].somModel.sram_ptr[1][24]=2;
sos_loop[0].somModel.sram_dat[1][25][0]=96'h699932;
sos_loop[0].somModel.sram_ptr[1][25]=2;
sos_loop[0].somModel.sram_dat[1][26][0]=96'h3c1356;
sos_loop[0].somModel.sram_ptr[1][26]=2;
sos_loop[0].somModel.sram_dat[1][27][0]=96'hda35e5;
sos_loop[0].somModel.sram_ptr[1][27]=2;
sos_loop[0].somModel.sram_dat[1][28][0]=96'hab08c2;
sos_loop[0].somModel.sram_ptr[1][28]=2;
sos_loop[0].somModel.sram_dat[1][29][0]=96'h55162c;
sos_loop[0].somModel.sram_ptr[1][29]=2;
sos_loop[0].somModel.sram_dat[1][30][0]=96'h48ac99;
sos_loop[0].somModel.sram_ptr[1][30]=2;
sos_loop[0].somModel.sram_dat[1][31][0]=96'hcf2b64;
sos_loop[0].somModel.sram_ptr[1][31]=2;
sos_loop[0].somModel.sram_dat[1][32][0]=96'he09d8f;
sos_loop[0].somModel.sram_ptr[1][32]=2;
sos_loop[0].somModel.sram_dat[1][33][0]=96'h1d11e0;
sos_loop[0].somModel.sram_ptr[1][33]=2;
sos_loop[0].somModel.sram_dat[1][34][0]=96'hdc6d6f;
sos_loop[0].somModel.sram_ptr[1][34]=2;
sos_loop[0].somModel.sram_dat[1][35][0]=96'h51d87e;
sos_loop[0].somModel.sram_ptr[1][35]=2;
sos_loop[0].somModel.sram_dat[1][36][0]=96'ha23c19;
sos_loop[0].somModel.sram_ptr[1][36]=2;
sos_loop[0].somModel.sram_dat[1][37][0]=96'ha8d569;
sos_loop[0].somModel.sram_ptr[1][37]=2;
sos_loop[0].somModel.sram_dat[1][38][0]=96'h9d9ed7;
sos_loop[0].somModel.sram_ptr[1][38]=2;
sos_loop[0].somModel.sram_dat[1][39][0]=96'h40e4d5;
sos_loop[0].somModel.sram_ptr[1][39]=2;
sos_loop[0].somModel.sram_dat[1][40][0]=96'h6b550f;
sos_loop[0].somModel.sram_ptr[1][40]=2;
sos_loop[0].somModel.sram_dat[1][41][0]=96'hb29e2e;
sos_loop[0].somModel.sram_ptr[1][41]=2;
sos_loop[0].somModel.sram_dat[1][42][0]=96'h2e7cf1;
sos_loop[0].somModel.sram_ptr[1][42]=2;
sos_loop[0].somModel.sram_dat[1][43][0]=96'h9200e3;
sos_loop[0].somModel.sram_ptr[1][43]=2;
sos_loop[0].somModel.sram_dat[1][44][0]=96'hd9b933;
sos_loop[0].somModel.sram_ptr[1][44]=2;
sos_loop[0].somModel.sram_dat[1][45][0]=96'hed726f;
sos_loop[0].somModel.sram_ptr[1][45]=2;
sos_loop[0].somModel.sram_dat[1][46][0]=96'h5a968d;
sos_loop[0].somModel.sram_ptr[1][46]=2;
sos_loop[0].somModel.sram_dat[1][47][0]=96'haa89df;
sos_loop[0].somModel.sram_ptr[1][47]=2;
sos_loop[0].somModel.sram_dat[1][48][0]=96'hc1a0ac;
sos_loop[0].somModel.sram_ptr[1][48]=2;
sos_loop[0].somModel.sram_dat[1][49][0]=96'h281727;
sos_loop[0].somModel.sram_ptr[1][49]=2;
sos_loop[0].somModel.sram_dat[1][50][0]=96'hfe964b;
sos_loop[0].somModel.sram_ptr[1][50]=2;
sos_loop[0].somModel.sram_dat[1][51][0]=96'h649d6a;
sos_loop[0].somModel.sram_ptr[1][51]=2;
sos_loop[0].somModel.sram_dat[1][52][0]=96'hb66d0f;
sos_loop[0].somModel.sram_ptr[1][52]=2;
sos_loop[0].somModel.sram_dat[1][53][0]=96'ha77176;
sos_loop[0].somModel.sram_ptr[1][53]=2;
sos_loop[0].somModel.sram_dat[1][54][0]=96'hab9e57;
sos_loop[0].somModel.sram_ptr[1][54]=2;
sos_loop[0].somModel.sram_dat[1][55][0]=96'he15190;
sos_loop[0].somModel.sram_ptr[1][55]=2;
sos_loop[0].somModel.sram_dat[1][56][0]=96'h935b3f;
sos_loop[0].somModel.sram_ptr[1][56]=2;
sos_loop[0].somModel.sram_dat[1][57][0]=96'h7d3e7;
sos_loop[0].somModel.sram_ptr[1][57]=2;
sos_loop[0].somModel.sram_dat[1][58][0]=96'hd866b3;
sos_loop[0].somModel.sram_ptr[1][58]=2;
sos_loop[0].somModel.sram_dat[1][59][0]=96'h4d2d96;
sos_loop[0].somModel.sram_ptr[1][59]=2;
sos_loop[0].somModel.sram_dat[1][60][0]=96'h932137;
sos_loop[0].somModel.sram_ptr[1][60]=2;
sos_loop[0].somModel.sram_dat[1][61][0]=96'hd76cda;
sos_loop[0].somModel.sram_ptr[1][61]=2;
sos_loop[0].somModel.sram_dat[1][62][0]=96'hcfb810;
sos_loop[0].somModel.sram_ptr[1][62]=2;
sos_loop[0].somModel.sram_dat[1][63][0]=96'h1f5e6f;
sos_loop[0].somModel.sram_ptr[1][63]=2;
sos_loop[0].somModel.sram_dat[1][64][0]=96'h866e5;
sos_loop[0].somModel.sram_ptr[1][64]=2;
sos_loop[0].somModel.sram_dat[1][65][0]=96'h552409;
sos_loop[0].somModel.sram_ptr[1][65]=2;
sos_loop[0].somModel.sram_dat[1][66][0]=96'h6819a;
sos_loop[0].somModel.sram_ptr[1][66]=2;
sos_loop[0].somModel.sram_dat[1][67][0]=96'hdabaa8;
sos_loop[0].somModel.sram_ptr[1][67]=2;
sos_loop[0].somModel.sram_dat[1][68][0]=96'h2fc8a9;
sos_loop[0].somModel.sram_ptr[1][68]=2;
sos_loop[0].somModel.sram_dat[1][69][0]=96'h5014e0;
sos_loop[0].somModel.sram_ptr[1][69]=2;
sos_loop[0].somModel.sram_dat[1][70][0]=96'hcc782f;
sos_loop[0].somModel.sram_ptr[1][70]=2;
sos_loop[0].somModel.sram_dat[1][71][0]=96'h6dae2a;
sos_loop[0].somModel.sram_ptr[1][71]=2;
sos_loop[0].somModel.sram_dat[1][72][0]=96'h39b496;
sos_loop[0].somModel.sram_ptr[1][72]=2;
sos_loop[0].somModel.sram_dat[1][73][0]=96'h1cae91;
sos_loop[0].somModel.sram_ptr[1][73]=2;
sos_loop[0].somModel.sram_dat[1][74][0]=96'hcaff50;
sos_loop[0].somModel.sram_ptr[1][74]=2;
sos_loop[0].somModel.sram_dat[1][75][0]=96'h33bd4;
sos_loop[0].somModel.sram_ptr[1][75]=2;
sos_loop[0].somModel.sram_dat[1][76][0]=96'h4cb006;
sos_loop[0].somModel.sram_ptr[1][76]=2;
sos_loop[0].somModel.sram_dat[1][77][0]=96'ha72599;
sos_loop[0].somModel.sram_ptr[1][77]=2;
sos_loop[0].somModel.sram_dat[1][78][0]=96'h19efb1;
sos_loop[0].somModel.sram_ptr[1][78]=2;
sos_loop[0].somModel.sram_dat[1][79][0]=96'hbc0688;
sos_loop[0].somModel.sram_ptr[1][79]=2;
sos_loop[0].somModel.sram_dat[1][80][0]=96'h37cb96;
sos_loop[0].somModel.sram_ptr[1][80]=2;
sos_loop[0].somModel.sram_dat[1][81][0]=96'h65d77e;
sos_loop[0].somModel.sram_ptr[1][81]=2;
sos_loop[0].somModel.sram_dat[1][82][0]=96'ha4e182;
sos_loop[0].somModel.sram_ptr[1][82]=2;
sos_loop[0].somModel.sram_dat[1][83][0]=96'hf9664b;
sos_loop[0].somModel.sram_ptr[1][83]=2;
sos_loop[0].somModel.sram_dat[1][84][0]=96'hd9d504;
sos_loop[0].somModel.sram_ptr[1][84]=2;
sos_loop[0].somModel.sram_dat[1][85][0]=96'hac6429;
sos_loop[0].somModel.sram_ptr[1][85]=2;
sos_loop[0].somModel.sram_dat[1][86][0]=96'h587b1;
sos_loop[0].somModel.sram_ptr[1][86]=2;
sos_loop[0].somModel.sram_dat[1][87][0]=96'h70b9ff;
sos_loop[0].somModel.sram_ptr[1][87]=2;
sos_loop[0].somModel.sram_dat[1][88][0]=96'h7817b3;
sos_loop[0].somModel.sram_ptr[1][88]=2;
sos_loop[0].somModel.sram_dat[1][89][0]=96'h5309c8;
sos_loop[0].somModel.sram_ptr[1][89]=2;
sos_loop[0].somModel.sram_dat[1][90][0]=96'h263667;
sos_loop[0].somModel.sram_ptr[1][90]=2;
sos_loop[0].somModel.sram_dat[1][91][0]=96'hbaef4d;
sos_loop[0].somModel.sram_ptr[1][91]=2;
sos_loop[0].somModel.sram_dat[1][92][0]=96'h9fe398;
sos_loop[0].somModel.sram_ptr[1][92]=2;
sos_loop[0].somModel.sram_dat[1][93][0]=96'hf404b2;
sos_loop[0].somModel.sram_ptr[1][93]=2;
sos_loop[0].somModel.sram_dat[1][94][0]=96'he66811;
sos_loop[0].somModel.sram_ptr[1][94]=2;
sos_loop[0].somModel.sram_dat[1][95][0]=96'h6c4854;
sos_loop[0].somModel.sram_ptr[1][95]=2;
sos_loop[0].somModel.sram_dat[1][96][0]=96'he41fbe;
sos_loop[0].somModel.sram_ptr[1][96]=2;
sos_loop[0].somModel.sram_dat[1][97][0]=96'hae926c;
sos_loop[0].somModel.sram_ptr[1][97]=2;
sos_loop[0].somModel.sram_dat[1][98][0]=96'h8b4995;
sos_loop[0].somModel.sram_ptr[1][98]=2;
sos_loop[0].somModel.sram_dat[1][99][0]=96'had9ee1;
sos_loop[0].somModel.sram_ptr[1][99]=2;
sos_loop[0].somModel.sram_dat[1][100][0]=96'he9cab6;
sos_loop[0].somModel.sram_ptr[1][100]=2;
sos_loop[0].somModel.sram_dat[1][101][0]=96'h190690;
sos_loop[0].somModel.sram_ptr[1][101]=2;
sos_loop[0].somModel.sram_dat[1][102][0]=96'h644cd1;
sos_loop[0].somModel.sram_ptr[1][102]=2;
sos_loop[0].somModel.sram_dat[1][103][0]=96'h193143;
sos_loop[0].somModel.sram_ptr[1][103]=2;
sos_loop[0].somModel.sram_dat[1][104][0]=96'hb38da9;
sos_loop[0].somModel.sram_ptr[1][104]=2;
sos_loop[0].somModel.sram_dat[1][105][0]=96'had42fb;
sos_loop[0].somModel.sram_ptr[1][105]=2;
sos_loop[0].somModel.sram_dat[1][106][0]=96'hf0c8e9;
sos_loop[0].somModel.sram_ptr[1][106]=2;
sos_loop[0].somModel.sram_dat[1][107][0]=96'hc63e22;
sos_loop[0].somModel.sram_ptr[1][107]=2;
sos_loop[0].somModel.sram_dat[1][108][0]=96'hceae4f;
sos_loop[0].somModel.sram_ptr[1][108]=2;
sos_loop[0].somModel.sram_dat[1][109][0]=96'h81fce1;
sos_loop[0].somModel.sram_ptr[1][109]=2;
sos_loop[0].somModel.sram_dat[1][110][0]=96'h6c8b8a;
sos_loop[0].somModel.sram_ptr[1][110]=2;
sos_loop[0].somModel.sram_dat[1][111][0]=96'hc9c607;
sos_loop[0].somModel.sram_ptr[1][111]=2;
sos_loop[0].somModel.sram_dat[1][112][0]=96'h84f36d;
sos_loop[0].somModel.sram_ptr[1][112]=2;
sos_loop[0].somModel.sram_dat[1][113][0]=96'h476c8a;
sos_loop[0].somModel.sram_ptr[1][113]=2;
sos_loop[0].somModel.sram_dat[1][114][0]=96'hd0a28d;
sos_loop[0].somModel.sram_ptr[1][114]=2;
sos_loop[0].somModel.sram_dat[1][115][0]=96'ha88374;
sos_loop[0].somModel.sram_ptr[1][115]=2;
sos_loop[0].somModel.sram_dat[1][116][0]=96'hec0149;
sos_loop[0].somModel.sram_ptr[1][116]=2;
sos_loop[0].somModel.sram_dat[1][117][0]=96'hd54c20;
sos_loop[0].somModel.sram_ptr[1][117]=2;
sos_loop[0].somModel.sram_dat[1][118][0]=96'h990140;
sos_loop[0].somModel.sram_ptr[1][118]=2;
sos_loop[0].somModel.sram_dat[1][119][0]=96'hd8c32b;
sos_loop[0].somModel.sram_ptr[1][119]=2;
sos_loop[0].somModel.sram_dat[1][120][0]=96'h9db7f1;
sos_loop[0].somModel.sram_ptr[1][120]=2;
sos_loop[0].somModel.sram_dat[1][121][0]=96'h4fa872;
sos_loop[0].somModel.sram_ptr[1][121]=2;
sos_loop[0].somModel.sram_dat[1][122][0]=96'hfa834c;
sos_loop[0].somModel.sram_ptr[1][122]=2;
sos_loop[0].somModel.sram_dat[1][123][0]=96'h640129;
sos_loop[0].somModel.sram_ptr[1][123]=2;
sos_loop[0].somModel.sram_dat[1][124][0]=96'h472ab0;
sos_loop[0].somModel.sram_ptr[1][124]=2;
sos_loop[0].somModel.sram_dat[1][125][0]=96'hde8fce;
sos_loop[0].somModel.sram_ptr[1][125]=2;
sos_loop[0].somModel.sram_dat[1][126][0]=96'he5dd77;
sos_loop[0].somModel.sram_ptr[1][126]=2;
sos_loop[0].somModel.sram_dat[1][127][0]=96'he2e528;
sos_loop[0].somModel.sram_ptr[1][127]=2;
sos_loop[0].somModel.sram_dat[1][128][0]=96'hc4a88f;
sos_loop[0].somModel.sram_ptr[1][128]=2;
sos_loop[0].somModel.sram_dat[1][129][0]=96'h36d132;
sos_loop[0].somModel.sram_ptr[1][129]=2;
sos_loop[0].somModel.sram_dat[1][130][0]=96'h103330;
sos_loop[0].somModel.sram_ptr[1][130]=2;
sos_loop[0].somModel.sram_dat[1][131][0]=96'h210b4b;
sos_loop[0].somModel.sram_ptr[1][131]=2;
sos_loop[0].somModel.sram_dat[1][132][0]=96'h23a29c;
sos_loop[0].somModel.sram_ptr[1][132]=2;
sos_loop[0].somModel.sram_dat[1][133][0]=96'h18d134;
sos_loop[0].somModel.sram_ptr[1][133]=2;
sos_loop[0].somModel.sram_dat[1][134][0]=96'h902d86;
sos_loop[0].somModel.sram_ptr[1][134]=2;
sos_loop[0].somModel.sram_dat[1][135][0]=96'h599e1e;
sos_loop[0].somModel.sram_ptr[1][135]=2;
sos_loop[0].somModel.sram_dat[1][136][0]=96'h8b80f3;
sos_loop[0].somModel.sram_ptr[1][136]=2;
sos_loop[0].somModel.sram_dat[1][137][0]=96'hfdd6d9;
sos_loop[0].somModel.sram_ptr[1][137]=2;
sos_loop[0].somModel.sram_dat[1][138][0]=96'ha822ed;
sos_loop[0].somModel.sram_ptr[1][138]=2;
sos_loop[0].somModel.sram_dat[1][139][0]=96'h325c6b;
sos_loop[0].somModel.sram_ptr[1][139]=2;
sos_loop[0].somModel.sram_dat[1][140][0]=96'hf3a0f1;
sos_loop[0].somModel.sram_ptr[1][140]=2;
sos_loop[0].somModel.sram_dat[1][141][0]=96'h40625f;
sos_loop[0].somModel.sram_ptr[1][141]=2;
sos_loop[0].somModel.sram_dat[1][142][0]=96'h62576;
sos_loop[0].somModel.sram_ptr[1][142]=2;
sos_loop[0].somModel.sram_dat[1][143][0]=96'h247741;
sos_loop[0].somModel.sram_ptr[1][143]=2;
sos_loop[0].somModel.sram_dat[1][144][0]=96'he66076;
sos_loop[0].somModel.sram_ptr[1][144]=2;
sos_loop[0].somModel.sram_dat[1][145][0]=96'ha1bfdb;
sos_loop[0].somModel.sram_ptr[1][145]=2;
sos_loop[0].somModel.sram_dat[1][146][0]=96'h733a59;
sos_loop[0].somModel.sram_ptr[1][146]=2;
sos_loop[0].somModel.sram_dat[1][147][0]=96'hd5364d;
sos_loop[0].somModel.sram_ptr[1][147]=2;
sos_loop[0].somModel.sram_dat[1][148][0]=96'hbf32c7;
sos_loop[0].somModel.sram_ptr[1][148]=2;
sos_loop[0].somModel.sram_dat[1][149][0]=96'hdc5dbf;
sos_loop[0].somModel.sram_ptr[1][149]=2;
sos_loop[0].somModel.sram_dat[1][150][0]=96'h9a93fb;
sos_loop[0].somModel.sram_ptr[1][150]=2;
sos_loop[0].somModel.sram_dat[1][151][0]=96'hcf1ba8;
sos_loop[0].somModel.sram_ptr[1][151]=2;
sos_loop[0].somModel.sram_dat[1][152][0]=96'h2a29f0;
sos_loop[0].somModel.sram_ptr[1][152]=2;
sos_loop[0].somModel.sram_dat[1][153][0]=96'hdbde8b;
sos_loop[0].somModel.sram_ptr[1][153]=2;
sos_loop[0].somModel.sram_dat[1][154][0]=96'h9fe4;
sos_loop[0].somModel.sram_ptr[1][154]=2;
sos_loop[0].somModel.sram_dat[1][155][0]=96'h180c0a;
sos_loop[0].somModel.sram_ptr[1][155]=2;
sos_loop[0].somModel.sram_dat[1][156][0]=96'h88f835;
sos_loop[0].somModel.sram_ptr[1][156]=2;
sos_loop[0].somModel.sram_dat[1][157][0]=96'h17109f;
sos_loop[0].somModel.sram_ptr[1][157]=2;
sos_loop[0].somModel.sram_dat[1][158][0]=96'h889713;
sos_loop[0].somModel.sram_ptr[1][158]=2;
sos_loop[0].somModel.sram_dat[1][159][0]=96'h41b6b6;
sos_loop[0].somModel.sram_ptr[1][159]=2;
sos_loop[0].somModel.sram_dat[1][160][0]=96'h864de9;
sos_loop[0].somModel.sram_ptr[1][160]=2;
sos_loop[0].somModel.sram_dat[1][161][0]=96'h7abce;
sos_loop[0].somModel.sram_ptr[1][161]=2;
sos_loop[0].somModel.sram_dat[1][162][0]=96'he12c35;
sos_loop[0].somModel.sram_ptr[1][162]=2;
sos_loop[0].somModel.sram_dat[1][163][0]=96'h301447;
sos_loop[0].somModel.sram_ptr[1][163]=2;
sos_loop[0].somModel.sram_dat[1][164][0]=96'h76b32;
sos_loop[0].somModel.sram_ptr[1][164]=2;
sos_loop[0].somModel.sram_dat[1][165][0]=96'h4b21b3;
sos_loop[0].somModel.sram_ptr[1][165]=2;
sos_loop[0].somModel.sram_dat[1][166][0]=96'ha87adb;
sos_loop[0].somModel.sram_ptr[1][166]=2;
sos_loop[0].somModel.sram_dat[1][167][0]=96'h8e26bd;
sos_loop[0].somModel.sram_ptr[1][167]=2;
sos_loop[0].somModel.sram_dat[1][168][0]=96'he69464;
sos_loop[0].somModel.sram_ptr[1][168]=2;
sos_loop[0].somModel.sram_dat[1][169][0]=96'hf1ae69;
sos_loop[0].somModel.sram_ptr[1][169]=2;
sos_loop[0].somModel.sram_dat[1][170][0]=96'h3aec7a;
sos_loop[0].somModel.sram_ptr[1][170]=2;
sos_loop[0].somModel.sram_dat[1][171][0]=96'hee62e2;
sos_loop[0].somModel.sram_ptr[1][171]=2;
sos_loop[0].somModel.sram_dat[1][172][0]=96'he8bc68;
sos_loop[0].somModel.sram_ptr[1][172]=2;
sos_loop[0].somModel.sram_dat[1][173][0]=96'h5b86a9;
sos_loop[0].somModel.sram_ptr[1][173]=2;
sos_loop[0].somModel.sram_dat[1][174][0]=96'h7871a5;
sos_loop[0].somModel.sram_ptr[1][174]=2;
sos_loop[0].somModel.sram_dat[1][175][0]=96'h55f1d9;
sos_loop[0].somModel.sram_ptr[1][175]=2;
sos_loop[0].somModel.sram_dat[1][176][0]=96'h96e694;
sos_loop[0].somModel.sram_ptr[1][176]=2;
sos_loop[0].somModel.sram_dat[1][177][0]=96'h1fe63b;
sos_loop[0].somModel.sram_ptr[1][177]=2;
sos_loop[0].somModel.sram_dat[1][178][0]=96'h806547;
sos_loop[0].somModel.sram_ptr[1][178]=2;
sos_loop[0].somModel.sram_dat[1][179][0]=96'h25c72f;
sos_loop[0].somModel.sram_ptr[1][179]=2;
sos_loop[0].somModel.sram_dat[1][180][0]=96'ha62af6;
sos_loop[0].somModel.sram_ptr[1][180]=2;
sos_loop[0].somModel.sram_dat[1][181][0]=96'h9d5417;
sos_loop[0].somModel.sram_ptr[1][181]=2;
sos_loop[0].somModel.sram_dat[1][182][0]=96'h2c51af;
sos_loop[0].somModel.sram_ptr[1][182]=2;
sos_loop[0].somModel.sram_dat[1][183][0]=96'h2f7ca4;
sos_loop[0].somModel.sram_ptr[1][183]=2;
sos_loop[0].somModel.sram_dat[1][184][0]=96'hc3d2cf;
sos_loop[0].somModel.sram_ptr[1][184]=2;
sos_loop[0].somModel.sram_dat[1][185][0]=96'h2f8d88;
sos_loop[0].somModel.sram_ptr[1][185]=2;
sos_loop[0].somModel.sram_dat[1][186][0]=96'h128302;
sos_loop[0].somModel.sram_ptr[1][186]=2;
sos_loop[0].somModel.sram_dat[1][187][0]=96'h3cc6e7;
sos_loop[0].somModel.sram_ptr[1][187]=2;
sos_loop[0].somModel.sram_dat[1][188][0]=96'hbebdfb;
sos_loop[0].somModel.sram_ptr[1][188]=2;
sos_loop[0].somModel.sram_dat[1][189][0]=96'haaacbb;
sos_loop[0].somModel.sram_ptr[1][189]=2;
sos_loop[0].somModel.sram_dat[1][190][0]=96'h35afca;
sos_loop[0].somModel.sram_ptr[1][190]=2;
sos_loop[0].somModel.sram_dat[1][191][0]=96'h3f635d;
sos_loop[0].somModel.sram_ptr[1][191]=2;
sos_loop[0].somModel.sram_dat[1][192][0]=96'h9dc27f;
sos_loop[0].somModel.sram_ptr[1][192]=2;
sos_loop[0].somModel.sram_dat[1][193][0]=96'hf64438;
sos_loop[0].somModel.sram_ptr[1][193]=2;
sos_loop[0].somModel.sram_dat[1][194][0]=96'h1cde19;
sos_loop[0].somModel.sram_ptr[1][194]=2;
sos_loop[0].somModel.sram_dat[1][195][0]=96'had0b70;
sos_loop[0].somModel.sram_ptr[1][195]=2;
sos_loop[0].somModel.sram_dat[1][196][0]=96'hb2a22c;
sos_loop[0].somModel.sram_ptr[1][196]=2;
sos_loop[0].somModel.sram_dat[1][197][0]=96'hc40815;
sos_loop[0].somModel.sram_ptr[1][197]=2;
sos_loop[0].somModel.sram_dat[1][198][0]=96'ha08a15;
sos_loop[0].somModel.sram_ptr[1][198]=2;
sos_loop[0].somModel.sram_dat[1][199][0]=96'h294352;
sos_loop[0].somModel.sram_ptr[1][199]=2;
sos_loop[0].somModel.sram_dat[1][200][0]=96'h9f922;
sos_loop[0].somModel.sram_ptr[1][200]=2;
sos_loop[0].somModel.sram_dat[1][201][0]=96'hc44933;
sos_loop[0].somModel.sram_ptr[1][201]=2;
sos_loop[0].somModel.sram_dat[1][202][0]=96'hcba9fb;
sos_loop[0].somModel.sram_ptr[1][202]=2;
sos_loop[0].somModel.sram_dat[1][203][0]=96'hcee397;
sos_loop[0].somModel.sram_ptr[1][203]=2;
sos_loop[0].somModel.sram_dat[1][204][0]=96'h5ab855;
sos_loop[0].somModel.sram_ptr[1][204]=2;
sos_loop[0].somModel.sram_dat[1][205][0]=96'hc37cff;
sos_loop[0].somModel.sram_ptr[1][205]=2;
sos_loop[0].somModel.sram_dat[1][206][0]=96'hf1815;
sos_loop[0].somModel.sram_ptr[1][206]=2;
sos_loop[0].somModel.sram_dat[1][207][0]=96'h1fecf8;
sos_loop[0].somModel.sram_ptr[1][207]=2;
sos_loop[0].somModel.sram_dat[1][208][0]=96'h2f0cd3;
sos_loop[0].somModel.sram_ptr[1][208]=2;
sos_loop[0].somModel.sram_dat[1][209][0]=96'hcdfdc7;
sos_loop[0].somModel.sram_ptr[1][209]=2;
sos_loop[0].somModel.sram_dat[1][210][0]=96'heada3f;
sos_loop[0].somModel.sram_ptr[1][210]=2;
sos_loop[0].somModel.sram_dat[1][211][0]=96'hc5239f;
sos_loop[0].somModel.sram_ptr[1][211]=2;
sos_loop[0].somModel.sram_dat[1][212][0]=96'h2e0306;
sos_loop[0].somModel.sram_ptr[1][212]=2;
sos_loop[0].somModel.sram_dat[1][213][0]=96'h9b50e8;
sos_loop[0].somModel.sram_ptr[1][213]=2;
sos_loop[0].somModel.sram_dat[1][214][0]=96'h244d2d;
sos_loop[0].somModel.sram_ptr[1][214]=2;
sos_loop[0].somModel.sram_dat[1][215][0]=96'hd04cf1;
sos_loop[0].somModel.sram_ptr[1][215]=2;
sos_loop[0].somModel.sram_dat[1][216][0]=96'h12056a;
sos_loop[0].somModel.sram_ptr[1][216]=2;
sos_loop[0].somModel.sram_dat[1][217][0]=96'h17ca62;
sos_loop[0].somModel.sram_ptr[1][217]=2;
sos_loop[0].somModel.sram_dat[1][218][0]=96'h3f7a75;
sos_loop[0].somModel.sram_ptr[1][218]=2;
sos_loop[0].somModel.sram_dat[1][219][0]=96'h7a839f;
sos_loop[0].somModel.sram_ptr[1][219]=2;
sos_loop[0].somModel.sram_dat[1][220][0]=96'h488d5;
sos_loop[0].somModel.sram_ptr[1][220]=2;
sos_loop[0].somModel.sram_dat[1][221][0]=96'h34ae81;
sos_loop[0].somModel.sram_ptr[1][221]=2;
sos_loop[0].somModel.sram_dat[1][222][0]=96'h1ee202;
sos_loop[0].somModel.sram_ptr[1][222]=2;
sos_loop[0].somModel.sram_dat[1][223][0]=96'h183ea5;
sos_loop[0].somModel.sram_ptr[1][223]=2;
sos_loop[0].somModel.sram_dat[1][224][0]=96'hc5cf43;
sos_loop[0].somModel.sram_ptr[1][224]=2;
sos_loop[0].somModel.sram_dat[1][225][0]=96'he2bc13;
sos_loop[0].somModel.sram_ptr[1][225]=2;
sos_loop[0].somModel.sram_dat[1][226][0]=96'h1fd051;
sos_loop[0].somModel.sram_ptr[1][226]=2;
sos_loop[0].somModel.sram_dat[1][227][0]=96'h1d970f;
sos_loop[0].somModel.sram_ptr[1][227]=2;
sos_loop[0].somModel.sram_dat[1][228][0]=96'hc403c7;
sos_loop[0].somModel.sram_ptr[1][228]=2;
sos_loop[0].somModel.sram_dat[1][229][0]=96'h88f8af;
sos_loop[0].somModel.sram_ptr[1][229]=2;
sos_loop[0].somModel.sram_dat[1][230][0]=96'h522f39;
sos_loop[0].somModel.sram_ptr[1][230]=2;
sos_loop[0].somModel.sram_dat[1][231][0]=96'hf385d1;
sos_loop[0].somModel.sram_ptr[1][231]=2;
sos_loop[0].somModel.sram_dat[1][232][0]=96'h9777c8;
sos_loop[0].somModel.sram_ptr[1][232]=2;
sos_loop[0].somModel.sram_dat[1][233][0]=96'hffee98;
sos_loop[0].somModel.sram_ptr[1][233]=2;
sos_loop[0].somModel.sram_dat[1][234][0]=96'h8f8852;
sos_loop[0].somModel.sram_ptr[1][234]=2;
sos_loop[0].somModel.sram_dat[1][235][0]=96'h22a823;
sos_loop[0].somModel.sram_ptr[1][235]=2;
sos_loop[0].somModel.sram_dat[1][236][0]=96'haabbdd;
sos_loop[0].somModel.sram_ptr[1][236]=2;
sos_loop[0].somModel.sram_dat[1][237][0]=96'hc4d792;
sos_loop[0].somModel.sram_ptr[1][237]=2;
sos_loop[0].somModel.sram_dat[1][238][0]=96'h1af82d;
sos_loop[0].somModel.sram_ptr[1][238]=2;
sos_loop[0].somModel.sram_dat[1][239][0]=96'h12e62a;
sos_loop[0].somModel.sram_ptr[1][239]=2;
sos_loop[0].somModel.sram_dat[1][240][0]=96'h84feb8;
sos_loop[0].somModel.sram_ptr[1][240]=2;
sos_loop[0].somModel.sram_dat[1][241][0]=96'he90935;
sos_loop[0].somModel.sram_ptr[1][241]=2;
sos_loop[0].somModel.sram_dat[1][242][0]=96'hdaeacf;
sos_loop[0].somModel.sram_ptr[1][242]=2;
sos_loop[0].somModel.sram_dat[1][243][0]=96'hf7fb36;
sos_loop[0].somModel.sram_ptr[1][243]=2;
sos_loop[0].somModel.sram_dat[1][244][0]=96'hb754c;
sos_loop[0].somModel.sram_ptr[1][244]=2;
sos_loop[0].somModel.sram_dat[1][245][0]=96'h72a0d2;
sos_loop[0].somModel.sram_ptr[1][245]=2;
sos_loop[0].somModel.sram_dat[1][246][0]=96'h14c7a8;
sos_loop[0].somModel.sram_ptr[1][246]=2;
sos_loop[0].somModel.sram_dat[1][247][0]=96'h2e7ccb;
sos_loop[0].somModel.sram_ptr[1][247]=2;
sos_loop[0].somModel.sram_dat[1][248][0]=96'h172d6b;
sos_loop[0].somModel.sram_ptr[1][248]=2;
sos_loop[0].somModel.sram_dat[1][249][0]=96'h5cbd69;
sos_loop[0].somModel.sram_ptr[1][249]=2;
sos_loop[0].somModel.sram_dat[1][250][0]=96'h838848;
sos_loop[0].somModel.sram_ptr[1][250]=2;
sos_loop[0].somModel.sram_dat[1][251][0]=96'he57f48;
sos_loop[0].somModel.sram_ptr[1][251]=2;
sos_loop[0].somModel.sram_dat[1][252][0]=96'h879954;
sos_loop[0].somModel.sram_ptr[1][252]=2;
sos_loop[0].somModel.sram_dat[1][253][0]=96'h3f3b48;
sos_loop[0].somModel.sram_ptr[1][253]=2;
sos_loop[0].somModel.sram_dat[1][254][0]=96'haa15a1;
sos_loop[0].somModel.sram_ptr[1][254]=2;
sos_loop[0].somModel.sram_dat[1][255][0]=96'h72e889;
sos_loop[0].somModel.sram_ptr[1][255]=2;
sos_loop[0].somModel.sram_dat[1][256][0]=96'h1b542;
sos_loop[0].somModel.sram_ptr[1][256]=2;
sos_loop[0].somModel.sram_dat[1][257][0]=96'h296632;
sos_loop[0].somModel.sram_ptr[1][257]=2;
sos_loop[0].somModel.sram_dat[1][258][0]=96'h38ad9e;
sos_loop[0].somModel.sram_ptr[1][258]=2;
sos_loop[0].somModel.sram_dat[1][259][0]=96'hdd5b20;
sos_loop[0].somModel.sram_ptr[1][259]=2;
sos_loop[0].somModel.sram_dat[1][260][0]=96'h7e3d3f;
sos_loop[0].somModel.sram_ptr[1][260]=2;
sos_loop[0].somModel.sram_dat[1][261][0]=96'hde577e;
sos_loop[0].somModel.sram_ptr[1][261]=2;
sos_loop[0].somModel.sram_dat[1][262][0]=96'h5f90c0;
sos_loop[0].somModel.sram_ptr[1][262]=2;
sos_loop[0].somModel.sram_dat[1][263][0]=96'hd30cb2;
sos_loop[0].somModel.sram_ptr[1][263]=2;
sos_loop[0].somModel.sram_dat[1][264][0]=96'h8ebe76;
sos_loop[0].somModel.sram_ptr[1][264]=2;
sos_loop[0].somModel.sram_dat[1][265][0]=96'h2d1e33;
sos_loop[0].somModel.sram_ptr[1][265]=2;
sos_loop[0].somModel.sram_dat[1][266][0]=96'h78e2fd;
sos_loop[0].somModel.sram_ptr[1][266]=2;
sos_loop[0].somModel.sram_dat[1][267][0]=96'h8595a0;
sos_loop[0].somModel.sram_ptr[1][267]=2;
sos_loop[0].somModel.sram_dat[1][268][0]=96'h4d7b60;
sos_loop[0].somModel.sram_ptr[1][268]=2;
sos_loop[0].somModel.sram_dat[1][269][0]=96'ha5d4d;
sos_loop[0].somModel.sram_ptr[1][269]=2;
sos_loop[0].somModel.sram_dat[1][270][0]=96'hb6a7b0;
sos_loop[0].somModel.sram_ptr[1][270]=2;
sos_loop[0].somModel.sram_dat[1][271][0]=96'hb9d0d8;
sos_loop[0].somModel.sram_ptr[1][271]=2;
sos_loop[0].somModel.sram_dat[1][272][0]=96'h7c54d0;
sos_loop[0].somModel.sram_ptr[1][272]=2;
sos_loop[0].somModel.sram_dat[1][273][0]=96'hfab;
sos_loop[0].somModel.sram_ptr[1][273]=2;
sos_loop[0].somModel.sram_dat[1][274][0]=96'h526452;
sos_loop[0].somModel.sram_ptr[1][274]=2;
sos_loop[0].somModel.sram_dat[1][275][0]=96'heea715;
sos_loop[0].somModel.sram_ptr[1][275]=2;
sos_loop[0].somModel.sram_dat[1][276][0]=96'hb958bc;
sos_loop[0].somModel.sram_ptr[1][276]=2;
sos_loop[0].somModel.sram_dat[1][277][0]=96'ha9b50c;
sos_loop[0].somModel.sram_ptr[1][277]=2;
sos_loop[0].somModel.sram_dat[1][278][0]=96'hfcbf5c;
sos_loop[0].somModel.sram_ptr[1][278]=2;
sos_loop[0].somModel.sram_dat[1][279][0]=96'hd7128e;
sos_loop[0].somModel.sram_ptr[1][279]=2;
sos_loop[0].somModel.sram_dat[1][280][0]=96'h287b14;
sos_loop[0].somModel.sram_ptr[1][280]=2;
sos_loop[0].somModel.sram_dat[1][281][0]=96'h99d893;
sos_loop[0].somModel.sram_ptr[1][281]=2;
sos_loop[0].somModel.sram_dat[1][282][0]=96'hce1be7;
sos_loop[0].somModel.sram_ptr[1][282]=2;
sos_loop[0].somModel.sram_dat[1][283][0]=96'h275c14;
sos_loop[0].somModel.sram_ptr[1][283]=2;
sos_loop[0].somModel.sram_dat[1][284][0]=96'hb2ecf6;
sos_loop[0].somModel.sram_ptr[1][284]=2;
sos_loop[0].somModel.sram_dat[1][285][0]=96'h32209f;
sos_loop[0].somModel.sram_ptr[1][285]=2;
sos_loop[0].somModel.sram_dat[1][286][0]=96'h8890e9;
sos_loop[0].somModel.sram_ptr[1][286]=2;
sos_loop[0].somModel.sram_dat[1][287][0]=96'h5df3a2;
sos_loop[0].somModel.sram_ptr[1][287]=2;
sos_loop[0].somModel.sram_dat[1][288][0]=96'h681f7e;
sos_loop[0].somModel.sram_ptr[1][288]=2;
sos_loop[0].somModel.sram_dat[1][289][0]=96'h52ac42;
sos_loop[0].somModel.sram_ptr[1][289]=2;
sos_loop[0].somModel.sram_dat[1][290][0]=96'h62b76d;
sos_loop[0].somModel.sram_ptr[1][290]=2;
sos_loop[0].somModel.sram_dat[1][291][0]=96'h2a3054;
sos_loop[0].somModel.sram_ptr[1][291]=2;
sos_loop[0].somModel.sram_dat[1][292][0]=96'ha6aacb;
sos_loop[0].somModel.sram_ptr[1][292]=2;
sos_loop[0].somModel.sram_dat[1][293][0]=96'hfad7b0;
sos_loop[0].somModel.sram_ptr[1][293]=2;
sos_loop[0].somModel.sram_dat[1][294][0]=96'he45af7;
sos_loop[0].somModel.sram_ptr[1][294]=2;
sos_loop[0].somModel.sram_dat[1][295][0]=96'h1b8312;
sos_loop[0].somModel.sram_ptr[1][295]=2;
sos_loop[0].somModel.sram_dat[1][296][0]=96'h4d7686;
sos_loop[0].somModel.sram_ptr[1][296]=2;
sos_loop[0].somModel.sram_dat[1][297][0]=96'h9e9f11;
sos_loop[0].somModel.sram_ptr[1][297]=2;
sos_loop[0].somModel.sram_dat[1][298][0]=96'h3752b8;
sos_loop[0].somModel.sram_ptr[1][298]=2;
sos_loop[0].somModel.sram_dat[1][299][0]=96'h9fff19;
sos_loop[0].somModel.sram_ptr[1][299]=2;
sos_loop[0].somModel.sram_dat[1][300][0]=96'h3deeb0;
sos_loop[0].somModel.sram_ptr[1][300]=2;
sos_loop[0].somModel.sram_dat[1][301][0]=96'h4d0cc0;
sos_loop[0].somModel.sram_ptr[1][301]=2;
sos_loop[0].somModel.sram_dat[1][302][0]=96'had4e0b;
sos_loop[0].somModel.sram_ptr[1][302]=2;
sos_loop[0].somModel.sram_dat[1][303][0]=96'hd93c76;
sos_loop[0].somModel.sram_ptr[1][303]=2;
sos_loop[0].somModel.sram_dat[1][304][0]=96'ha363f3;
sos_loop[0].somModel.sram_ptr[1][304]=2;
sos_loop[0].somModel.sram_dat[1][305][0]=96'hfe7a4a;
sos_loop[0].somModel.sram_ptr[1][305]=2;
sos_loop[0].somModel.sram_dat[1][306][0]=96'h6750fd;
sos_loop[0].somModel.sram_ptr[1][306]=2;
sos_loop[0].somModel.sram_dat[1][307][0]=96'hfa4199;
sos_loop[0].somModel.sram_ptr[1][307]=2;
sos_loop[0].somModel.sram_dat[1][308][0]=96'hd91f85;
sos_loop[0].somModel.sram_ptr[1][308]=2;
sos_loop[0].somModel.sram_dat[1][309][0]=96'h6021c5;
sos_loop[0].somModel.sram_ptr[1][309]=2;
sos_loop[0].somModel.sram_dat[1][310][0]=96'hb7fc65;
sos_loop[0].somModel.sram_ptr[1][310]=2;
sos_loop[0].somModel.sram_dat[1][311][0]=96'hd6e41;
sos_loop[0].somModel.sram_ptr[1][311]=2;
sos_loop[0].somModel.sram_dat[1][312][0]=96'h1fc6a1;
sos_loop[0].somModel.sram_ptr[1][312]=2;
sos_loop[0].somModel.sram_dat[1][313][0]=96'hd152b0;
sos_loop[0].somModel.sram_ptr[1][313]=2;
sos_loop[0].somModel.sram_dat[1][314][0]=96'h2f8780;
sos_loop[0].somModel.sram_ptr[1][314]=2;
sos_loop[0].somModel.sram_dat[1][315][0]=96'ha9948;
sos_loop[0].somModel.sram_ptr[1][315]=2;
sos_loop[0].somModel.sram_dat[1][316][0]=96'h249ab8;
sos_loop[0].somModel.sram_ptr[1][316]=2;
sos_loop[0].somModel.sram_dat[1][317][0]=96'h472875;
sos_loop[0].somModel.sram_ptr[1][317]=2;
sos_loop[0].somModel.sram_dat[1][318][0]=96'h6d2196;
sos_loop[0].somModel.sram_ptr[1][318]=2;
sos_loop[0].somModel.sram_dat[1][319][0]=96'h10373f;
sos_loop[0].somModel.sram_ptr[1][319]=2;
sos_loop[0].somModel.sram_dat[1][320][0]=96'hc0f50e;
sos_loop[0].somModel.sram_ptr[1][320]=2;
sos_loop[0].somModel.sram_dat[1][321][0]=96'hdd84a8;
sos_loop[0].somModel.sram_ptr[1][321]=2;
sos_loop[0].somModel.sram_dat[1][322][0]=96'h324444;
sos_loop[0].somModel.sram_ptr[1][322]=2;
sos_loop[0].somModel.sram_dat[1][323][0]=96'hb11fe3;
sos_loop[0].somModel.sram_ptr[1][323]=2;
sos_loop[0].somModel.sram_dat[1][324][0]=96'hd3c003;
sos_loop[0].somModel.sram_ptr[1][324]=2;
sos_loop[0].somModel.sram_dat[1][325][0]=96'h22c068;
sos_loop[0].somModel.sram_ptr[1][325]=2;
sos_loop[0].somModel.sram_dat[1][326][0]=96'h200557;
sos_loop[0].somModel.sram_ptr[1][326]=2;
sos_loop[0].somModel.sram_dat[1][327][0]=96'hd760d5;
sos_loop[0].somModel.sram_ptr[1][327]=2;
sos_loop[0].somModel.sram_dat[1][328][0]=96'h404d84;
sos_loop[0].somModel.sram_ptr[1][328]=2;
sos_loop[0].somModel.sram_dat[1][329][0]=96'h38a6a0;
sos_loop[0].somModel.sram_ptr[1][329]=2;
sos_loop[0].somModel.sram_dat[1][330][0]=96'h3a4640;
sos_loop[0].somModel.sram_ptr[1][330]=2;
sos_loop[0].somModel.sram_dat[1][331][0]=96'h4a10b1;
sos_loop[0].somModel.sram_ptr[1][331]=2;
sos_loop[0].somModel.sram_dat[1][332][0]=96'hb30115;
sos_loop[0].somModel.sram_ptr[1][332]=2;
sos_loop[0].somModel.sram_dat[1][333][0]=96'h8aeaa5;
sos_loop[0].somModel.sram_ptr[1][333]=2;
sos_loop[0].somModel.sram_dat[1][334][0]=96'hf1cc59;
sos_loop[0].somModel.sram_ptr[1][334]=2;
sos_loop[0].somModel.sram_dat[1][335][0]=96'h7f6f35;
sos_loop[0].somModel.sram_ptr[1][335]=2;
sos_loop[0].somModel.sram_dat[1][336][0]=96'h465838;
sos_loop[0].somModel.sram_ptr[1][336]=2;
sos_loop[0].somModel.sram_dat[1][337][0]=96'hc08db5;
sos_loop[0].somModel.sram_ptr[1][337]=2;
sos_loop[0].somModel.sram_dat[1][338][0]=96'hfd7be1;
sos_loop[0].somModel.sram_ptr[1][338]=2;
sos_loop[0].somModel.sram_dat[1][339][0]=96'ha0f3;
sos_loop[0].somModel.sram_ptr[1][339]=2;
sos_loop[0].somModel.sram_dat[1][340][0]=96'hb91869;
sos_loop[0].somModel.sram_ptr[1][340]=2;
sos_loop[0].somModel.sram_dat[1][341][0]=96'hc0ad63;
sos_loop[0].somModel.sram_ptr[1][341]=2;
sos_loop[0].somModel.sram_dat[1][342][0]=96'hb08e22;
sos_loop[0].somModel.sram_ptr[1][342]=2;
sos_loop[0].somModel.sram_dat[1][343][0]=96'hf68553;
sos_loop[0].somModel.sram_ptr[1][343]=2;
sos_loop[0].somModel.sram_dat[1][344][0]=96'h64927f;
sos_loop[0].somModel.sram_ptr[1][344]=2;
sos_loop[0].somModel.sram_dat[1][345][0]=96'h83a02e;
sos_loop[0].somModel.sram_ptr[1][345]=2;
sos_loop[0].somModel.sram_dat[1][346][0]=96'hbe5a96;
sos_loop[0].somModel.sram_ptr[1][346]=2;
sos_loop[0].somModel.sram_dat[1][347][0]=96'h6e40d1;
sos_loop[0].somModel.sram_ptr[1][347]=2;
sos_loop[0].somModel.sram_dat[1][348][0]=96'hf76daa;
sos_loop[0].somModel.sram_ptr[1][348]=2;
sos_loop[0].somModel.sram_dat[1][349][0]=96'h260806;
sos_loop[0].somModel.sram_ptr[1][349]=2;
sos_loop[0].somModel.sram_dat[1][350][0]=96'haaf348;
sos_loop[0].somModel.sram_ptr[1][350]=2;
sos_loop[0].somModel.sram_dat[1][351][0]=96'hbe1a7;
sos_loop[0].somModel.sram_ptr[1][351]=2;
sos_loop[0].somModel.sram_dat[1][352][0]=96'ha59283;
sos_loop[0].somModel.sram_ptr[1][352]=2;
sos_loop[0].somModel.sram_dat[1][353][0]=96'h9fd1ab;
sos_loop[0].somModel.sram_ptr[1][353]=2;
sos_loop[0].somModel.sram_dat[1][354][0]=96'h8acbff;
sos_loop[0].somModel.sram_ptr[1][354]=2;
sos_loop[0].somModel.sram_dat[1][355][0]=96'h4deca7;
sos_loop[0].somModel.sram_ptr[1][355]=2;
sos_loop[0].somModel.sram_dat[1][356][0]=96'h28e13a;
sos_loop[0].somModel.sram_ptr[1][356]=2;
sos_loop[0].somModel.sram_dat[1][357][0]=96'ha299ca;
sos_loop[0].somModel.sram_ptr[1][357]=2;
sos_loop[0].somModel.sram_dat[1][358][0]=96'h99a477;
sos_loop[0].somModel.sram_ptr[1][358]=2;
sos_loop[0].somModel.sram_dat[1][359][0]=96'h44a766;
sos_loop[0].somModel.sram_ptr[1][359]=2;
sos_loop[0].somModel.sram_dat[1][360][0]=96'hd3a394;
sos_loop[0].somModel.sram_ptr[1][360]=2;
sos_loop[0].somModel.sram_dat[1][361][0]=96'hecc3e8;
sos_loop[0].somModel.sram_ptr[1][361]=2;
sos_loop[0].somModel.sram_dat[1][362][0]=96'hebab0e;
sos_loop[0].somModel.sram_ptr[1][362]=2;
sos_loop[0].somModel.sram_dat[1][363][0]=96'h7f07a0;
sos_loop[0].somModel.sram_ptr[1][363]=2;
sos_loop[0].somModel.sram_dat[1][364][0]=96'h1940da;
sos_loop[0].somModel.sram_ptr[1][364]=2;
sos_loop[0].somModel.sram_dat[1][365][0]=96'hdd77fd;
sos_loop[0].somModel.sram_ptr[1][365]=2;
sos_loop[0].somModel.sram_dat[1][366][0]=96'h27a422;
sos_loop[0].somModel.sram_ptr[1][366]=2;
sos_loop[0].somModel.sram_dat[1][367][0]=96'he19559;
sos_loop[0].somModel.sram_ptr[1][367]=2;
sos_loop[0].somModel.sram_dat[1][368][0]=96'h8d63;
sos_loop[0].somModel.sram_ptr[1][368]=2;
sos_loop[0].somModel.sram_dat[1][369][0]=96'h1193c;
sos_loop[0].somModel.sram_ptr[1][369]=2;
sos_loop[0].somModel.sram_dat[1][370][0]=96'h46a7c0;
sos_loop[0].somModel.sram_ptr[1][370]=2;
sos_loop[0].somModel.sram_dat[1][371][0]=96'hc71745;
sos_loop[0].somModel.sram_ptr[1][371]=2;
sos_loop[0].somModel.sram_dat[1][372][0]=96'hee0321;
sos_loop[0].somModel.sram_ptr[1][372]=2;
sos_loop[0].somModel.sram_dat[1][373][0]=96'h21c943;
sos_loop[0].somModel.sram_ptr[1][373]=2;
sos_loop[0].somModel.sram_dat[1][374][0]=96'h5334c6;
sos_loop[0].somModel.sram_ptr[1][374]=2;
sos_loop[0].somModel.sram_dat[1][375][0]=96'hcbd414;
sos_loop[0].somModel.sram_ptr[1][375]=2;
sos_loop[0].somModel.sram_dat[1][376][0]=96'hab0538;
sos_loop[0].somModel.sram_ptr[1][376]=2;
sos_loop[0].somModel.sram_dat[1][377][0]=96'hf176c0;
sos_loop[0].somModel.sram_ptr[1][377]=2;
sos_loop[0].somModel.sram_dat[1][378][0]=96'h8512ed;
sos_loop[0].somModel.sram_ptr[1][378]=2;
sos_loop[0].somModel.sram_dat[1][379][0]=96'ha0128d;
sos_loop[0].somModel.sram_ptr[1][379]=2;
sos_loop[0].somModel.sram_dat[1][380][0]=96'hdb3124;
sos_loop[0].somModel.sram_ptr[1][380]=2;
sos_loop[0].somModel.sram_dat[1][381][0]=96'h3d7888;
sos_loop[0].somModel.sram_ptr[1][381]=2;
sos_loop[0].somModel.sram_dat[1][382][0]=96'h6f91b;
sos_loop[0].somModel.sram_ptr[1][382]=2;
sos_loop[0].somModel.sram_dat[1][383][0]=96'hb21e43;
sos_loop[0].somModel.sram_ptr[1][383]=2;
sos_loop[0].somModel.sram_dat[1][384][0]=96'h8de00c;
sos_loop[0].somModel.sram_ptr[1][384]=2;
sos_loop[0].somModel.sram_dat[1][385][0]=96'had6a91;
sos_loop[0].somModel.sram_ptr[1][385]=2;
sos_loop[0].somModel.sram_dat[1][386][0]=96'h9982b5;
sos_loop[0].somModel.sram_ptr[1][386]=2;
sos_loop[0].somModel.sram_dat[1][387][0]=96'hf936b6;
sos_loop[0].somModel.sram_ptr[1][387]=2;
sos_loop[0].somModel.sram_dat[1][388][0]=96'hfb8434;
sos_loop[0].somModel.sram_ptr[1][388]=2;
sos_loop[0].somModel.sram_dat[1][389][0]=96'h61ac31;
sos_loop[0].somModel.sram_ptr[1][389]=2;
sos_loop[0].somModel.sram_dat[1][390][0]=96'hd66;
sos_loop[0].somModel.sram_ptr[1][390]=2;
sos_loop[0].somModel.sram_dat[1][391][0]=96'hcb4d6b;
sos_loop[0].somModel.sram_ptr[1][391]=2;
sos_loop[0].somModel.sram_dat[1][392][0]=96'h952555;
sos_loop[0].somModel.sram_ptr[1][392]=2;
sos_loop[0].somModel.sram_dat[1][393][0]=96'hd662de;
sos_loop[0].somModel.sram_ptr[1][393]=2;
sos_loop[0].somModel.sram_dat[1][394][0]=96'haa0ea6;
sos_loop[0].somModel.sram_ptr[1][394]=2;
sos_loop[0].somModel.sram_dat[1][395][0]=96'hba2e0f;
sos_loop[0].somModel.sram_ptr[1][395]=2;
sos_loop[0].somModel.sram_dat[1][396][0]=96'hf7491c;
sos_loop[0].somModel.sram_ptr[1][396]=2;
sos_loop[0].somModel.sram_dat[1][397][0]=96'h8d68ee;
sos_loop[0].somModel.sram_ptr[1][397]=2;
sos_loop[0].somModel.sram_dat[1][398][0]=96'ha366a5;
sos_loop[0].somModel.sram_ptr[1][398]=2;
sos_loop[0].somModel.sram_dat[1][399][0]=96'h7672fe;
sos_loop[0].somModel.sram_ptr[1][399]=2;
sos_loop[0].somModel.sram_dat[1][400][0]=96'h4e0e5b;
sos_loop[0].somModel.sram_ptr[1][400]=2;
sos_loop[0].somModel.sram_dat[1][401][0]=96'hf69f93;
sos_loop[0].somModel.sram_ptr[1][401]=2;
sos_loop[0].somModel.sram_dat[1][402][0]=96'hdc64a3;
sos_loop[0].somModel.sram_ptr[1][402]=2;
sos_loop[0].somModel.sram_dat[1][403][0]=96'h3e36d7;
sos_loop[0].somModel.sram_ptr[1][403]=2;
sos_loop[0].somModel.sram_dat[1][404][0]=96'h20cd14;
sos_loop[0].somModel.sram_ptr[1][404]=2;
sos_loop[0].somModel.sram_dat[1][405][0]=96'hfd80ee;
sos_loop[0].somModel.sram_ptr[1][405]=2;
sos_loop[0].somModel.sram_dat[1][406][0]=96'h14a853;
sos_loop[0].somModel.sram_ptr[1][406]=2;
sos_loop[0].somModel.sram_dat[1][407][0]=96'hd34e71;
sos_loop[0].somModel.sram_ptr[1][407]=2;
sos_loop[0].somModel.sram_dat[1][408][0]=96'h4da43e;
sos_loop[0].somModel.sram_ptr[1][408]=2;
sos_loop[0].somModel.sram_dat[1][409][0]=96'h2dcdd0;
sos_loop[0].somModel.sram_ptr[1][409]=2;
sos_loop[0].somModel.sram_dat[1][410][0]=96'hff51e4;
sos_loop[0].somModel.sram_ptr[1][410]=2;
sos_loop[0].somModel.sram_dat[1][411][0]=96'h5e4c3b;
sos_loop[0].somModel.sram_ptr[1][411]=2;
sos_loop[0].somModel.sram_dat[1][412][0]=96'h919a50;
sos_loop[0].somModel.sram_ptr[1][412]=2;
sos_loop[0].somModel.sram_dat[1][413][0]=96'h5c6f6;
sos_loop[0].somModel.sram_ptr[1][413]=2;
sos_loop[0].somModel.sram_dat[1][414][0]=96'h4880e1;
sos_loop[0].somModel.sram_ptr[1][414]=2;
sos_loop[0].somModel.sram_dat[1][415][0]=96'hb52f6e;
sos_loop[0].somModel.sram_ptr[1][415]=2;
sos_loop[0].somModel.sram_dat[1][416][0]=96'h6330f5;
sos_loop[0].somModel.sram_ptr[1][416]=2;
sos_loop[0].somModel.sram_dat[1][417][0]=96'h87589c;
sos_loop[0].somModel.sram_ptr[1][417]=2;
sos_loop[0].somModel.sram_dat[1][418][0]=96'hae87c5;
sos_loop[0].somModel.sram_ptr[1][418]=2;
sos_loop[0].somModel.sram_dat[1][419][0]=96'h88b591;
sos_loop[0].somModel.sram_ptr[1][419]=2;
sos_loop[0].somModel.sram_dat[1][420][0]=96'ha9681c;
sos_loop[0].somModel.sram_ptr[1][420]=2;
sos_loop[0].somModel.sram_dat[1][421][0]=96'h5bfe8c;
sos_loop[0].somModel.sram_ptr[1][421]=2;
sos_loop[0].somModel.sram_dat[1][422][0]=96'hfeeabb;
sos_loop[0].somModel.sram_ptr[1][422]=2;
sos_loop[0].somModel.sram_dat[1][423][0]=96'h5bfef3;
sos_loop[0].somModel.sram_ptr[1][423]=2;
sos_loop[0].somModel.sram_dat[1][424][0]=96'hc439f5;
sos_loop[0].somModel.sram_ptr[1][424]=2;
sos_loop[0].somModel.sram_dat[1][425][0]=96'hcbb611;
sos_loop[0].somModel.sram_ptr[1][425]=2;
sos_loop[0].somModel.sram_dat[1][426][0]=96'h6bf841;
sos_loop[0].somModel.sram_ptr[1][426]=2;
sos_loop[0].somModel.sram_dat[1][427][0]=96'h14eb96;
sos_loop[0].somModel.sram_ptr[1][427]=2;
sos_loop[0].somModel.sram_dat[1][428][0]=96'hcb6ce3;
sos_loop[0].somModel.sram_ptr[1][428]=2;
sos_loop[0].somModel.sram_dat[1][429][0]=96'hbe0907;
sos_loop[0].somModel.sram_ptr[1][429]=2;
sos_loop[0].somModel.sram_dat[1][430][0]=96'hf515b5;
sos_loop[0].somModel.sram_ptr[1][430]=2;
sos_loop[0].somModel.sram_dat[1][431][0]=96'hd4b21b;
sos_loop[0].somModel.sram_ptr[1][431]=2;
sos_loop[0].somModel.sram_dat[1][432][0]=96'haed1b5;
sos_loop[0].somModel.sram_ptr[1][432]=2;
sos_loop[0].somModel.sram_dat[1][433][0]=96'h187e1;
sos_loop[0].somModel.sram_ptr[1][433]=2;
sos_loop[0].somModel.sram_dat[1][434][0]=96'h3bf896;
sos_loop[0].somModel.sram_ptr[1][434]=2;
sos_loop[0].somModel.sram_dat[1][435][0]=96'hd53055;
sos_loop[0].somModel.sram_ptr[1][435]=2;
sos_loop[0].somModel.sram_dat[1][436][0]=96'hd85a46;
sos_loop[0].somModel.sram_ptr[1][436]=2;
sos_loop[0].somModel.sram_dat[1][437][0]=96'hb70da5;
sos_loop[0].somModel.sram_ptr[1][437]=2;
sos_loop[0].somModel.sram_dat[1][438][0]=96'hf14efb;
sos_loop[0].somModel.sram_ptr[1][438]=2;
sos_loop[0].somModel.sram_dat[1][439][0]=96'hceed54;
sos_loop[0].somModel.sram_ptr[1][439]=2;
sos_loop[0].somModel.sram_dat[1][440][0]=96'h1c63cc;
sos_loop[0].somModel.sram_ptr[1][440]=2;
sos_loop[0].somModel.sram_dat[1][441][0]=96'h2e657b;
sos_loop[0].somModel.sram_ptr[1][441]=2;
sos_loop[0].somModel.sram_dat[1][442][0]=96'h1b7bb1;
sos_loop[0].somModel.sram_ptr[1][442]=2;
sos_loop[0].somModel.sram_dat[1][443][0]=96'ha490bb;
sos_loop[0].somModel.sram_ptr[1][443]=2;
sos_loop[0].somModel.sram_dat[1][444][0]=96'h77f7c3;
sos_loop[0].somModel.sram_ptr[1][444]=2;
sos_loop[0].somModel.sram_dat[1][445][0]=96'hce3879;
sos_loop[0].somModel.sram_ptr[1][445]=2;
sos_loop[0].somModel.sram_dat[1][446][0]=96'h3d62f7;
sos_loop[0].somModel.sram_ptr[1][446]=2;
sos_loop[0].somModel.sram_dat[1][447][0]=96'hd3c317;
sos_loop[0].somModel.sram_ptr[1][447]=2;
sos_loop[0].somModel.sram_dat[1][448][0]=96'hcd4052;
sos_loop[0].somModel.sram_ptr[1][448]=2;
sos_loop[0].somModel.sram_dat[1][449][0]=96'h366029;
sos_loop[0].somModel.sram_ptr[1][449]=2;
sos_loop[0].somModel.sram_dat[1][450][0]=96'h249c31;
sos_loop[0].somModel.sram_ptr[1][450]=2;
sos_loop[0].somModel.sram_dat[1][451][0]=96'hf85353;
sos_loop[0].somModel.sram_ptr[1][451]=2;
sos_loop[0].somModel.sram_dat[1][452][0]=96'hba861d;
sos_loop[0].somModel.sram_ptr[1][452]=2;
sos_loop[0].somModel.sram_dat[1][453][0]=96'h7b4f14;
sos_loop[0].somModel.sram_ptr[1][453]=2;
sos_loop[0].somModel.sram_dat[1][454][0]=96'he9a8b0;
sos_loop[0].somModel.sram_ptr[1][454]=2;
sos_loop[0].somModel.sram_dat[1][455][0]=96'h48daff;
sos_loop[0].somModel.sram_ptr[1][455]=2;
sos_loop[0].somModel.sram_dat[1][456][0]=96'h9eeb3;
sos_loop[0].somModel.sram_ptr[1][456]=2;
sos_loop[0].somModel.sram_dat[1][457][0]=96'h1ea67;
sos_loop[0].somModel.sram_ptr[1][457]=2;
sos_loop[0].somModel.sram_dat[1][458][0]=96'hb2c532;
sos_loop[0].somModel.sram_ptr[1][458]=2;
sos_loop[0].somModel.sram_dat[1][459][0]=96'h8cdabd;
sos_loop[0].somModel.sram_ptr[1][459]=2;
sos_loop[0].somModel.sram_dat[1][460][0]=96'he33611;
sos_loop[0].somModel.sram_ptr[1][460]=2;
sos_loop[0].somModel.sram_dat[1][461][0]=96'h888646;
sos_loop[0].somModel.sram_ptr[1][461]=2;
sos_loop[0].somModel.sram_dat[1][462][0]=96'h7532ec;
sos_loop[0].somModel.sram_ptr[1][462]=2;
sos_loop[0].somModel.sram_dat[1][463][0]=96'hef77eb;
sos_loop[0].somModel.sram_ptr[1][463]=2;
sos_loop[0].somModel.sram_dat[1][464][0]=96'h836a74;
sos_loop[0].somModel.sram_ptr[1][464]=2;
sos_loop[0].somModel.sram_dat[1][465][0]=96'h60abde;
sos_loop[0].somModel.sram_ptr[1][465]=2;
sos_loop[0].somModel.sram_dat[1][466][0]=96'h1fb207;
sos_loop[0].somModel.sram_ptr[1][466]=2;
sos_loop[0].somModel.sram_dat[1][467][0]=96'h1fd4bb;
sos_loop[0].somModel.sram_ptr[1][467]=2;
sos_loop[0].somModel.sram_dat[1][468][0]=96'he37673;
sos_loop[0].somModel.sram_ptr[1][468]=2;
sos_loop[0].somModel.sram_dat[1][469][0]=96'he78f3e;
sos_loop[0].somModel.sram_ptr[1][469]=2;
sos_loop[0].somModel.sram_dat[1][470][0]=96'hf089bc;
sos_loop[0].somModel.sram_ptr[1][470]=2;
sos_loop[0].somModel.sram_dat[1][471][0]=96'h989a46;
sos_loop[0].somModel.sram_ptr[1][471]=2;
sos_loop[0].somModel.sram_dat[1][472][0]=96'h4872d;
sos_loop[0].somModel.sram_ptr[1][472]=2;
sos_loop[0].somModel.sram_dat[1][473][0]=96'h7d4a59;
sos_loop[0].somModel.sram_ptr[1][473]=2;
sos_loop[0].somModel.sram_dat[1][474][0]=96'h79148c;
sos_loop[0].somModel.sram_ptr[1][474]=2;
sos_loop[0].somModel.sram_dat[1][475][0]=96'hca4d53;
sos_loop[0].somModel.sram_ptr[1][475]=2;
sos_loop[0].somModel.sram_dat[1][476][0]=96'h318859;
sos_loop[0].somModel.sram_ptr[1][476]=2;
sos_loop[0].somModel.sram_dat[1][477][0]=96'hd19af7;
sos_loop[0].somModel.sram_ptr[1][477]=2;
sos_loop[0].somModel.sram_dat[1][478][0]=96'h270545;
sos_loop[0].somModel.sram_ptr[1][478]=2;
sos_loop[0].somModel.sram_dat[1][479][0]=96'h94a8f5;
sos_loop[0].somModel.sram_ptr[1][479]=2;
sos_loop[0].somModel.sram_dat[1][480][0]=96'hfd4a65;
sos_loop[0].somModel.sram_ptr[1][480]=2;
sos_loop[0].somModel.sram_dat[1][481][0]=96'h14a4ed;
sos_loop[0].somModel.sram_ptr[1][481]=2;
sos_loop[0].somModel.sram_dat[1][482][0]=96'hb279ba;
sos_loop[0].somModel.sram_ptr[1][482]=2;
sos_loop[0].somModel.sram_dat[1][483][0]=96'h63905b;
sos_loop[0].somModel.sram_ptr[1][483]=2;
sos_loop[0].somModel.sram_dat[1][484][0]=96'h528285;
sos_loop[0].somModel.sram_ptr[1][484]=2;
sos_loop[0].somModel.sram_dat[1][485][0]=96'hbd6eb1;
sos_loop[0].somModel.sram_ptr[1][485]=2;
sos_loop[0].somModel.sram_dat[1][486][0]=96'h136e6c;
sos_loop[0].somModel.sram_ptr[1][486]=2;
sos_loop[0].somModel.sram_dat[1][487][0]=96'h9b3456;
sos_loop[0].somModel.sram_ptr[1][487]=2;
sos_loop[0].somModel.sram_dat[1][488][0]=96'h254c0a;
sos_loop[0].somModel.sram_ptr[1][488]=2;
sos_loop[0].somModel.sram_dat[1][489][0]=96'hec438c;
sos_loop[0].somModel.sram_ptr[1][489]=2;
sos_loop[0].somModel.sram_dat[1][490][0]=96'h84699d;
sos_loop[0].somModel.sram_ptr[1][490]=2;
sos_loop[0].somModel.sram_dat[1][491][0]=96'hd0224;
sos_loop[0].somModel.sram_ptr[1][491]=2;
sos_loop[0].somModel.sram_dat[1][492][0]=96'hc49916;
sos_loop[0].somModel.sram_ptr[1][492]=2;
sos_loop[0].somModel.sram_dat[1][493][0]=96'hff4173;
sos_loop[0].somModel.sram_ptr[1][493]=2;
sos_loop[0].somModel.sram_dat[1][494][0]=96'h81bccf;
sos_loop[0].somModel.sram_ptr[1][494]=2;
sos_loop[0].somModel.sram_dat[1][495][0]=96'h6fed17;
sos_loop[0].somModel.sram_ptr[1][495]=2;
sos_loop[0].somModel.sram_dat[1][496][0]=96'h2329d9;
sos_loop[0].somModel.sram_ptr[1][496]=2;
sos_loop[0].somModel.sram_dat[1][497][0]=96'he35295;
sos_loop[0].somModel.sram_ptr[1][497]=2;
sos_loop[0].somModel.sram_dat[1][498][0]=96'h97a6ce;
sos_loop[0].somModel.sram_ptr[1][498]=2;
sos_loop[0].somModel.sram_dat[1][499][0]=96'h7355fd;
sos_loop[0].somModel.sram_ptr[1][499]=2;
sos_loop[0].somModel.sram_dat[1][500][0]=96'hb5e794;
sos_loop[0].somModel.sram_ptr[1][500]=2;
sos_loop[0].somModel.sram_dat[1][501][0]=96'h3295ab;
sos_loop[0].somModel.sram_ptr[1][501]=2;
sos_loop[0].somModel.sram_dat[1][502][0]=96'heca5ce;
sos_loop[0].somModel.sram_ptr[1][502]=2;
sos_loop[0].somModel.sram_dat[1][503][0]=96'h87bf14;
sos_loop[0].somModel.sram_ptr[1][503]=2;
sos_loop[0].somModel.sram_dat[1][504][0]=96'ha166f5;
sos_loop[0].somModel.sram_ptr[1][504]=2;
sos_loop[0].somModel.sram_dat[1][505][0]=96'hc0b98a;
sos_loop[0].somModel.sram_ptr[1][505]=2;
sos_loop[0].somModel.sram_dat[1][506][0]=96'h452cdc;
sos_loop[0].somModel.sram_ptr[1][506]=2;
sos_loop[0].somModel.sram_dat[1][507][0]=96'h78e1e0;
sos_loop[0].somModel.sram_ptr[1][507]=2;
sos_loop[0].somModel.sram_dat[1][508][0]=96'h92eb8c;
sos_loop[0].somModel.sram_ptr[1][508]=2;
sos_loop[0].somModel.sram_dat[1][509][0]=96'h129629;
sos_loop[0].somModel.sram_ptr[1][509]=2;
sos_loop[0].somModel.sram_dat[1][510][0]=96'hbc837b;
sos_loop[0].somModel.sram_ptr[1][510]=2;
sos_loop[0].somModel.sram_dat[1][511][0]=96'h9cda8f;
sos_loop[0].somModel.sram_ptr[1][511]=2;
sos_loop[0].somModel.sram_dat[1][512][0]=96'h3e36f7;
sos_loop[0].somModel.sram_ptr[1][512]=2;
sos_loop[0].somModel.sram_dat[1][513][0]=96'h8a27cd;
sos_loop[0].somModel.sram_ptr[1][513]=2;
sos_loop[0].somModel.sram_dat[1][514][0]=96'h462c62;
sos_loop[0].somModel.sram_ptr[1][514]=2;
sos_loop[0].somModel.sram_dat[1][515][0]=96'hdfcade;
sos_loop[0].somModel.sram_ptr[1][515]=2;
sos_loop[0].somModel.sram_dat[1][516][0]=96'h8989c8;
sos_loop[0].somModel.sram_ptr[1][516]=2;
sos_loop[0].somModel.sram_dat[1][517][0]=96'h6c0294;
sos_loop[0].somModel.sram_ptr[1][517]=2;
sos_loop[0].somModel.sram_dat[1][518][0]=96'hbcd2eb;
sos_loop[0].somModel.sram_ptr[1][518]=2;
sos_loop[0].somModel.sram_dat[1][519][0]=96'h3bff68;
sos_loop[0].somModel.sram_ptr[1][519]=2;
sos_loop[0].somModel.sram_dat[1][520][0]=96'h6b9b27;
sos_loop[0].somModel.sram_ptr[1][520]=2;
sos_loop[0].somModel.sram_dat[1][521][0]=96'h22b3ea;
sos_loop[0].somModel.sram_ptr[1][521]=2;
sos_loop[0].somModel.sram_dat[1][522][0]=96'h41688a;
sos_loop[0].somModel.sram_ptr[1][522]=2;
sos_loop[0].somModel.sram_dat[1][523][0]=96'he21345;
sos_loop[0].somModel.sram_ptr[1][523]=2;
sos_loop[0].somModel.sram_dat[1][524][0]=96'h73d32b;
sos_loop[0].somModel.sram_ptr[1][524]=2;
sos_loop[0].somModel.sram_dat[1][525][0]=96'ha2a953;
sos_loop[0].somModel.sram_ptr[1][525]=2;
sos_loop[0].somModel.sram_dat[1][526][0]=96'h4e430c;
sos_loop[0].somModel.sram_ptr[1][526]=2;
sos_loop[0].somModel.sram_dat[1][527][0]=96'h64d84c;
sos_loop[0].somModel.sram_ptr[1][527]=2;
sos_loop[0].somModel.sram_dat[1][528][0]=96'h2f0b4c;
sos_loop[0].somModel.sram_ptr[1][528]=2;
sos_loop[0].somModel.sram_dat[1][529][0]=96'h3b69f1;
sos_loop[0].somModel.sram_ptr[1][529]=2;
sos_loop[0].somModel.sram_dat[1][530][0]=96'hac0c0;
sos_loop[0].somModel.sram_ptr[1][530]=2;
sos_loop[0].somModel.sram_dat[1][531][0]=96'h2cb8c;
sos_loop[0].somModel.sram_ptr[1][531]=2;
sos_loop[0].somModel.sram_dat[1][532][0]=96'hc8973d;
sos_loop[0].somModel.sram_ptr[1][532]=2;
sos_loop[0].somModel.sram_dat[1][533][0]=96'h63403b;
sos_loop[0].somModel.sram_ptr[1][533]=2;
sos_loop[0].somModel.sram_dat[1][534][0]=96'h3b10ba;
sos_loop[0].somModel.sram_ptr[1][534]=2;
sos_loop[0].somModel.sram_dat[1][535][0]=96'h2ce7ba;
sos_loop[0].somModel.sram_ptr[1][535]=2;
sos_loop[0].somModel.sram_dat[1][536][0]=96'hea87;
sos_loop[0].somModel.sram_ptr[1][536]=2;
sos_loop[0].somModel.sram_dat[1][537][0]=96'h50badf;
sos_loop[0].somModel.sram_ptr[1][537]=2;
sos_loop[0].somModel.sram_dat[1][538][0]=96'h5b2fbb;
sos_loop[0].somModel.sram_ptr[1][538]=2;
sos_loop[0].somModel.sram_dat[1][539][0]=96'hac32d9;
sos_loop[0].somModel.sram_ptr[1][539]=2;
sos_loop[0].somModel.sram_dat[1][540][0]=96'h175207;
sos_loop[0].somModel.sram_ptr[1][540]=2;
sos_loop[0].somModel.sram_dat[1][541][0]=96'hce27f9;
sos_loop[0].somModel.sram_ptr[1][541]=2;
sos_loop[0].somModel.sram_dat[1][542][0]=96'h75d740;
sos_loop[0].somModel.sram_ptr[1][542]=2;
sos_loop[0].somModel.sram_dat[1][543][0]=96'h76d79a;
sos_loop[0].somModel.sram_ptr[1][543]=2;
sos_loop[0].somModel.sram_dat[1][544][0]=96'h7390f8;
sos_loop[0].somModel.sram_ptr[1][544]=2;
sos_loop[0].somModel.sram_dat[1][545][0]=96'hb963bf;
sos_loop[0].somModel.sram_ptr[1][545]=2;
sos_loop[0].somModel.sram_dat[1][546][0]=96'h26405;
sos_loop[0].somModel.sram_ptr[1][546]=2;
sos_loop[0].somModel.sram_dat[1][547][0]=96'ha04b21;
sos_loop[0].somModel.sram_ptr[1][547]=2;
sos_loop[0].somModel.sram_dat[1][548][0]=96'ha30541;
sos_loop[0].somModel.sram_ptr[1][548]=2;
sos_loop[0].somModel.sram_dat[1][549][0]=96'h8927b6;
sos_loop[0].somModel.sram_ptr[1][549]=2;
sos_loop[0].somModel.sram_dat[1][550][0]=96'h9cc1c0;
sos_loop[0].somModel.sram_ptr[1][550]=2;
sos_loop[0].somModel.sram_dat[1][551][0]=96'h3ba3f5;
sos_loop[0].somModel.sram_ptr[1][551]=2;
sos_loop[0].somModel.sram_dat[1][552][0]=96'h352e1d;
sos_loop[0].somModel.sram_ptr[1][552]=2;
sos_loop[0].somModel.sram_dat[1][553][0]=96'hc2fbc1;
sos_loop[0].somModel.sram_ptr[1][553]=2;
sos_loop[0].somModel.sram_dat[1][554][0]=96'h4cbb09;
sos_loop[0].somModel.sram_ptr[1][554]=2;
sos_loop[0].somModel.sram_dat[1][555][0]=96'hffbbbf;
sos_loop[0].somModel.sram_ptr[1][555]=2;
sos_loop[0].somModel.sram_dat[1][556][0]=96'hb682c8;
sos_loop[0].somModel.sram_ptr[1][556]=2;
sos_loop[0].somModel.sram_dat[1][557][0]=96'h52c4da;
sos_loop[0].somModel.sram_ptr[1][557]=2;
sos_loop[0].somModel.sram_dat[1][558][0]=96'h312a41;
sos_loop[0].somModel.sram_ptr[1][558]=2;
sos_loop[0].somModel.sram_dat[1][559][0]=96'h8b4d5;
sos_loop[0].somModel.sram_ptr[1][559]=2;
sos_loop[0].somModel.sram_dat[1][560][0]=96'hf3a2ad;
sos_loop[0].somModel.sram_ptr[1][560]=2;
sos_loop[0].somModel.sram_dat[1][561][0]=96'h6e7c4f;
sos_loop[0].somModel.sram_ptr[1][561]=2;
sos_loop[0].somModel.sram_dat[1][562][0]=96'hded8dc;
sos_loop[0].somModel.sram_ptr[1][562]=2;
sos_loop[0].somModel.sram_dat[1][563][0]=96'h1dc81;
sos_loop[0].somModel.sram_ptr[1][563]=2;
sos_loop[0].somModel.sram_dat[1][564][0]=96'hfbaf9;
sos_loop[0].somModel.sram_ptr[1][564]=2;
sos_loop[0].somModel.sram_dat[1][565][0]=96'h61584b;
sos_loop[0].somModel.sram_ptr[1][565]=2;
sos_loop[0].somModel.sram_dat[1][566][0]=96'h7649b8;
sos_loop[0].somModel.sram_ptr[1][566]=2;
sos_loop[0].somModel.sram_dat[1][567][0]=96'h5f5cd1;
sos_loop[0].somModel.sram_ptr[1][567]=2;
sos_loop[0].somModel.sram_dat[1][568][0]=96'hf10131;
sos_loop[0].somModel.sram_ptr[1][568]=2;
sos_loop[0].somModel.sram_dat[1][569][0]=96'h72671c;
sos_loop[0].somModel.sram_ptr[1][569]=2;
sos_loop[0].somModel.sram_dat[1][570][0]=96'hd3785d;
sos_loop[0].somModel.sram_ptr[1][570]=2;
sos_loop[0].somModel.sram_dat[1][571][0]=96'ha29593;
sos_loop[0].somModel.sram_ptr[1][571]=2;
sos_loop[0].somModel.sram_dat[1][572][0]=96'h954c60;
sos_loop[0].somModel.sram_ptr[1][572]=2;
sos_loop[0].somModel.sram_dat[1][573][0]=96'hc17e8e;
sos_loop[0].somModel.sram_ptr[1][573]=2;
sos_loop[0].somModel.sram_dat[1][574][0]=96'h9a7ba;
sos_loop[0].somModel.sram_ptr[1][574]=2;
sos_loop[0].somModel.sram_dat[1][575][0]=96'h7072f3;
sos_loop[0].somModel.sram_ptr[1][575]=2;
sos_loop[0].somModel.sram_dat[1][576][0]=96'h78fcbf;
sos_loop[0].somModel.sram_ptr[1][576]=2;
sos_loop[0].somModel.sram_dat[1][577][0]=96'h43c1b7;
sos_loop[0].somModel.sram_ptr[1][577]=2;
sos_loop[0].somModel.sram_dat[1][578][0]=96'hb08007;
sos_loop[0].somModel.sram_ptr[1][578]=2;
sos_loop[0].somModel.sram_dat[1][579][0]=96'h150566;
sos_loop[0].somModel.sram_ptr[1][579]=2;
sos_loop[0].somModel.sram_dat[1][580][0]=96'ha9a978;
sos_loop[0].somModel.sram_ptr[1][580]=2;
sos_loop[0].somModel.sram_dat[1][581][0]=96'hc86b86;
sos_loop[0].somModel.sram_ptr[1][581]=2;
sos_loop[0].somModel.sram_dat[1][582][0]=96'hf6a9b4;
sos_loop[0].somModel.sram_ptr[1][582]=2;
sos_loop[0].somModel.sram_dat[1][583][0]=96'hbd5e1d;
sos_loop[0].somModel.sram_ptr[1][583]=2;
sos_loop[0].somModel.sram_dat[1][584][0]=96'h6bdf3d;
sos_loop[0].somModel.sram_ptr[1][584]=2;
sos_loop[0].somModel.sram_dat[1][585][0]=96'h8848ec;
sos_loop[0].somModel.sram_ptr[1][585]=2;
sos_loop[0].somModel.sram_dat[1][586][0]=96'h2de4cb;
sos_loop[0].somModel.sram_ptr[1][586]=2;
sos_loop[0].somModel.sram_dat[1][587][0]=96'h729081;
sos_loop[0].somModel.sram_ptr[1][587]=2;
sos_loop[0].somModel.sram_dat[1][588][0]=96'h6a8d3d;
sos_loop[0].somModel.sram_ptr[1][588]=2;
sos_loop[0].somModel.sram_dat[1][589][0]=96'hb986e7;
sos_loop[0].somModel.sram_ptr[1][589]=2;
sos_loop[0].somModel.sram_dat[1][590][0]=96'h53a9dc;
sos_loop[0].somModel.sram_ptr[1][590]=2;
sos_loop[0].somModel.sram_dat[1][591][0]=96'h495aab;
sos_loop[0].somModel.sram_ptr[1][591]=2;
sos_loop[0].somModel.sram_dat[1][592][0]=96'h2243c5;
sos_loop[0].somModel.sram_ptr[1][592]=2;
sos_loop[0].somModel.sram_dat[1][593][0]=96'h932bc5;
sos_loop[0].somModel.sram_ptr[1][593]=2;
sos_loop[0].somModel.sram_dat[1][594][0]=96'hc7e5a1;
sos_loop[0].somModel.sram_ptr[1][594]=2;
sos_loop[0].somModel.sram_dat[1][595][0]=96'h519f51;
sos_loop[0].somModel.sram_ptr[1][595]=2;
sos_loop[0].somModel.sram_dat[1][596][0]=96'h31d9d3;
sos_loop[0].somModel.sram_ptr[1][596]=2;
sos_loop[0].somModel.sram_dat[1][597][0]=96'h6c648c;
sos_loop[0].somModel.sram_ptr[1][597]=2;
sos_loop[0].somModel.sram_dat[1][598][0]=96'hca4098;
sos_loop[0].somModel.sram_ptr[1][598]=2;
sos_loop[0].somModel.sram_dat[1][599][0]=96'he6aa63;
sos_loop[0].somModel.sram_ptr[1][599]=2;
sos_loop[0].somModel.sram_dat[1][600][0]=96'h9898d6;
sos_loop[0].somModel.sram_ptr[1][600]=2;
sos_loop[0].somModel.sram_dat[1][601][0]=96'h2e0ee6;
sos_loop[0].somModel.sram_ptr[1][601]=2;
sos_loop[0].somModel.sram_dat[1][602][0]=96'h7de959;
sos_loop[0].somModel.sram_ptr[1][602]=2;
sos_loop[0].somModel.sram_dat[1][603][0]=96'h22ed5e;
sos_loop[0].somModel.sram_ptr[1][603]=2;
sos_loop[0].somModel.sram_dat[1][604][0]=96'hef9cd4;
sos_loop[0].somModel.sram_ptr[1][604]=2;
sos_loop[0].somModel.sram_dat[1][605][0]=96'h9e573b;
sos_loop[0].somModel.sram_ptr[1][605]=2;
sos_loop[0].somModel.sram_dat[1][606][0]=96'ha4a6bf;
sos_loop[0].somModel.sram_ptr[1][606]=2;
sos_loop[0].somModel.sram_dat[1][607][0]=96'h96fae7;
sos_loop[0].somModel.sram_ptr[1][607]=2;
sos_loop[0].somModel.sram_dat[1][608][0]=96'hcdbaec;
sos_loop[0].somModel.sram_ptr[1][608]=2;
sos_loop[0].somModel.sram_dat[1][609][0]=96'hf9a463;
sos_loop[0].somModel.sram_ptr[1][609]=2;
sos_loop[0].somModel.sram_dat[1][610][0]=96'h4e36e0;
sos_loop[0].somModel.sram_ptr[1][610]=2;
sos_loop[0].somModel.sram_dat[1][611][0]=96'hf0a7a9;
sos_loop[0].somModel.sram_ptr[1][611]=2;
sos_loop[0].somModel.sram_dat[1][612][0]=96'h1ae7e7;
sos_loop[0].somModel.sram_ptr[1][612]=2;
sos_loop[0].somModel.sram_dat[1][613][0]=96'hfacdcc;
sos_loop[0].somModel.sram_ptr[1][613]=2;
sos_loop[0].somModel.sram_dat[1][614][0]=96'h57f90;
sos_loop[0].somModel.sram_ptr[1][614]=2;
sos_loop[0].somModel.sram_dat[1][615][0]=96'hb782da;
sos_loop[0].somModel.sram_ptr[1][615]=2;
sos_loop[0].somModel.sram_dat[1][616][0]=96'h68b3;
sos_loop[0].somModel.sram_ptr[1][616]=2;
sos_loop[0].somModel.sram_dat[1][617][0]=96'h3a8542;
sos_loop[0].somModel.sram_ptr[1][617]=2;
sos_loop[0].somModel.sram_dat[1][618][0]=96'h662a36;
sos_loop[0].somModel.sram_ptr[1][618]=2;
sos_loop[0].somModel.sram_dat[1][619][0]=96'hc447e7;
sos_loop[0].somModel.sram_ptr[1][619]=2;
sos_loop[0].somModel.sram_dat[1][620][0]=96'h428275;
sos_loop[0].somModel.sram_ptr[1][620]=2;
sos_loop[0].somModel.sram_dat[1][621][0]=96'h207e9f;
sos_loop[0].somModel.sram_ptr[1][621]=2;
sos_loop[0].somModel.sram_dat[1][622][0]=96'hb5de9b;
sos_loop[0].somModel.sram_ptr[1][622]=2;
sos_loop[0].somModel.sram_dat[1][623][0]=96'hbdfb18;
sos_loop[0].somModel.sram_ptr[1][623]=2;
sos_loop[0].somModel.sram_dat[1][624][0]=96'h3a7a85;
sos_loop[0].somModel.sram_ptr[1][624]=2;
sos_loop[0].somModel.sram_dat[1][625][0]=96'h6b085d;
sos_loop[0].somModel.sram_ptr[1][625]=2;
sos_loop[0].somModel.sram_dat[1][626][0]=96'he56816;
sos_loop[0].somModel.sram_ptr[1][626]=2;
sos_loop[0].somModel.sram_dat[1][627][0]=96'h18d22b;
sos_loop[0].somModel.sram_ptr[1][627]=2;
sos_loop[0].somModel.sram_dat[1][628][0]=96'hfd73c1;
sos_loop[0].somModel.sram_ptr[1][628]=2;
sos_loop[0].somModel.sram_dat[1][629][0]=96'hf65166;
sos_loop[0].somModel.sram_ptr[1][629]=2;
sos_loop[0].somModel.sram_dat[1][630][0]=96'haea4f6;
sos_loop[0].somModel.sram_ptr[1][630]=2;
sos_loop[0].somModel.sram_dat[1][631][0]=96'h378ad7;
sos_loop[0].somModel.sram_ptr[1][631]=2;
sos_loop[0].somModel.sram_dat[1][632][0]=96'h7215cb;
sos_loop[0].somModel.sram_ptr[1][632]=2;
sos_loop[0].somModel.sram_dat[1][633][0]=96'h4370d3;
sos_loop[0].somModel.sram_ptr[1][633]=2;
sos_loop[0].somModel.sram_dat[1][634][0]=96'he0bb48;
sos_loop[0].somModel.sram_ptr[1][634]=2;
sos_loop[0].somModel.sram_dat[1][635][0]=96'hdd2dbc;
sos_loop[0].somModel.sram_ptr[1][635]=2;
sos_loop[0].somModel.sram_dat[1][636][0]=96'hd10c0d;
sos_loop[0].somModel.sram_ptr[1][636]=2;
sos_loop[0].somModel.sram_dat[1][637][0]=96'h45ca7b;
sos_loop[0].somModel.sram_ptr[1][637]=2;
sos_loop[0].somModel.sram_dat[1][638][0]=96'h50ec64;
sos_loop[0].somModel.sram_ptr[1][638]=2;
sos_loop[0].somModel.sram_dat[1][639][0]=96'h906144;
sos_loop[0].somModel.sram_ptr[1][639]=2;
sos_loop[0].somModel.sram_dat[1][640][0]=96'h112dc1;
sos_loop[0].somModel.sram_ptr[1][640]=2;
sos_loop[0].somModel.sram_dat[1][641][0]=96'h5b36ae;
sos_loop[0].somModel.sram_ptr[1][641]=2;
sos_loop[0].somModel.sram_dat[1][642][0]=96'h6a5c37;
sos_loop[0].somModel.sram_ptr[1][642]=2;
sos_loop[0].somModel.sram_dat[1][643][0]=96'h24a942;
sos_loop[0].somModel.sram_ptr[1][643]=2;
sos_loop[0].somModel.sram_dat[1][644][0]=96'h48e2b;
sos_loop[0].somModel.sram_ptr[1][644]=2;
sos_loop[0].somModel.sram_dat[1][645][0]=96'h77fa27;
sos_loop[0].somModel.sram_ptr[1][645]=2;
sos_loop[0].somModel.sram_dat[1][646][0]=96'h78b151;
sos_loop[0].somModel.sram_ptr[1][646]=2;
sos_loop[0].somModel.sram_dat[1][647][0]=96'ha47604;
sos_loop[0].somModel.sram_ptr[1][647]=2;
sos_loop[0].somModel.sram_dat[1][648][0]=96'h594a3f;
sos_loop[0].somModel.sram_ptr[1][648]=2;
sos_loop[0].somModel.sram_dat[1][649][0]=96'haf2e91;
sos_loop[0].somModel.sram_ptr[1][649]=2;
sos_loop[0].somModel.sram_dat[1][650][0]=96'h54f406;
sos_loop[0].somModel.sram_ptr[1][650]=2;
sos_loop[0].somModel.sram_dat[1][651][0]=96'hdbd353;
sos_loop[0].somModel.sram_ptr[1][651]=2;
sos_loop[0].somModel.sram_dat[1][652][0]=96'ha961f7;
sos_loop[0].somModel.sram_ptr[1][652]=2;
sos_loop[0].somModel.sram_dat[1][653][0]=96'h655384;
sos_loop[0].somModel.sram_ptr[1][653]=2;
sos_loop[0].somModel.sram_dat[1][654][0]=96'h1b8b2;
sos_loop[0].somModel.sram_ptr[1][654]=2;
sos_loop[0].somModel.sram_dat[1][655][0]=96'hb646a0;
sos_loop[0].somModel.sram_ptr[1][655]=2;
sos_loop[0].somModel.sram_dat[1][656][0]=96'hc35541;
sos_loop[0].somModel.sram_ptr[1][656]=2;
sos_loop[0].somModel.sram_dat[1][657][0]=96'haa459d;
sos_loop[0].somModel.sram_ptr[1][657]=2;
sos_loop[0].somModel.sram_dat[1][658][0]=96'h759b4f;
sos_loop[0].somModel.sram_ptr[1][658]=2;
sos_loop[0].somModel.sram_dat[1][659][0]=96'h10b764;
sos_loop[0].somModel.sram_ptr[1][659]=2;
sos_loop[0].somModel.sram_dat[1][660][0]=96'h7f2ca2;
sos_loop[0].somModel.sram_ptr[1][660]=2;
sos_loop[0].somModel.sram_dat[1][661][0]=96'h9605;
sos_loop[0].somModel.sram_ptr[1][661]=2;
sos_loop[0].somModel.sram_dat[1][662][0]=96'h880ee7;
sos_loop[0].somModel.sram_ptr[1][662]=2;
sos_loop[0].somModel.sram_dat[1][663][0]=96'heced99;
sos_loop[0].somModel.sram_ptr[1][663]=2;
sos_loop[0].somModel.sram_dat[1][664][0]=96'h8a05ca;
sos_loop[0].somModel.sram_ptr[1][664]=2;
sos_loop[0].somModel.sram_dat[1][665][0]=96'h66baf9;
sos_loop[0].somModel.sram_ptr[1][665]=2;
sos_loop[0].somModel.sram_dat[1][666][0]=96'h96805d;
sos_loop[0].somModel.sram_ptr[1][666]=2;
sos_loop[0].somModel.sram_dat[1][667][0]=96'he3de2;
sos_loop[0].somModel.sram_ptr[1][667]=2;
sos_loop[0].somModel.sram_dat[1][668][0]=96'h15e3df;
sos_loop[0].somModel.sram_ptr[1][668]=2;
sos_loop[0].somModel.sram_dat[1][669][0]=96'ha47712;
sos_loop[0].somModel.sram_ptr[1][669]=2;
sos_loop[0].somModel.sram_dat[1][670][0]=96'h1932f3;
sos_loop[0].somModel.sram_ptr[1][670]=2;
sos_loop[0].somModel.sram_dat[1][671][0]=96'h15d54c;
sos_loop[0].somModel.sram_ptr[1][671]=2;
sos_loop[0].somModel.sram_dat[1][672][0]=96'h8e6097;
sos_loop[0].somModel.sram_ptr[1][672]=2;
sos_loop[0].somModel.sram_dat[1][673][0]=96'h26723;
sos_loop[0].somModel.sram_ptr[1][673]=2;
sos_loop[0].somModel.sram_dat[1][674][0]=96'h2d4201;
sos_loop[0].somModel.sram_ptr[1][674]=2;
sos_loop[0].somModel.sram_dat[1][675][0]=96'h64a019;
sos_loop[0].somModel.sram_ptr[1][675]=2;
sos_loop[0].somModel.sram_dat[1][676][0]=96'h52068;
sos_loop[0].somModel.sram_ptr[1][676]=2;
sos_loop[0].somModel.sram_dat[1][677][0]=96'h4fc87f;
sos_loop[0].somModel.sram_ptr[1][677]=2;
sos_loop[0].somModel.sram_dat[1][678][0]=96'h354c4a;
sos_loop[0].somModel.sram_ptr[1][678]=2;
sos_loop[0].somModel.sram_dat[1][679][0]=96'hc084df;
sos_loop[0].somModel.sram_ptr[1][679]=2;
sos_loop[0].somModel.sram_dat[1][680][0]=96'he3af6c;
sos_loop[0].somModel.sram_ptr[1][680]=2;
sos_loop[0].somModel.sram_dat[1][681][0]=96'h9b4c6a;
sos_loop[0].somModel.sram_ptr[1][681]=2;
sos_loop[0].somModel.sram_dat[1][682][0]=96'h4fe061;
sos_loop[0].somModel.sram_ptr[1][682]=2;
sos_loop[0].somModel.sram_dat[1][683][0]=96'h668b54;
sos_loop[0].somModel.sram_ptr[1][683]=2;
sos_loop[0].somModel.sram_dat[1][684][0]=96'hb7d2fa;
sos_loop[0].somModel.sram_ptr[1][684]=2;
sos_loop[0].somModel.sram_dat[1][685][0]=96'h7b394b;
sos_loop[0].somModel.sram_ptr[1][685]=2;
sos_loop[0].somModel.sram_dat[1][686][0]=96'ha0d693;
sos_loop[0].somModel.sram_ptr[1][686]=2;
sos_loop[0].somModel.sram_dat[1][687][0]=96'hecb9e8;
sos_loop[0].somModel.sram_ptr[1][687]=2;
sos_loop[0].somModel.sram_dat[1][688][0]=96'hfa6dcb;
sos_loop[0].somModel.sram_ptr[1][688]=2;
sos_loop[0].somModel.sram_dat[1][689][0]=96'h549727;
sos_loop[0].somModel.sram_ptr[1][689]=2;
sos_loop[0].somModel.sram_dat[1][690][0]=96'h563be7;
sos_loop[0].somModel.sram_ptr[1][690]=2;
sos_loop[0].somModel.sram_dat[1][691][0]=96'hefc0f2;
sos_loop[0].somModel.sram_ptr[1][691]=2;
sos_loop[0].somModel.sram_dat[1][692][0]=96'hc5e4f2;
sos_loop[0].somModel.sram_ptr[1][692]=2;
sos_loop[0].somModel.sram_dat[1][693][0]=96'h97e2e2;
sos_loop[0].somModel.sram_ptr[1][693]=2;
sos_loop[0].somModel.sram_dat[1][694][0]=96'hd71d42;
sos_loop[0].somModel.sram_ptr[1][694]=2;
sos_loop[0].somModel.sram_dat[1][695][0]=96'h2cc08f;
sos_loop[0].somModel.sram_ptr[1][695]=2;
sos_loop[0].somModel.sram_dat[1][696][0]=96'h6e18f9;
sos_loop[0].somModel.sram_ptr[1][696]=2;
sos_loop[0].somModel.sram_dat[1][697][0]=96'hfdf59;
sos_loop[0].somModel.sram_ptr[1][697]=2;
sos_loop[0].somModel.sram_dat[1][698][0]=96'h8f22b0;
sos_loop[0].somModel.sram_ptr[1][698]=2;
sos_loop[0].somModel.sram_dat[1][699][0]=96'hf70e50;
sos_loop[0].somModel.sram_ptr[1][699]=2;
sos_loop[0].somModel.sram_dat[1][700][0]=96'h65c364;
sos_loop[0].somModel.sram_ptr[1][700]=2;
sos_loop[0].somModel.cfg_tbl_sel[1] = 1;
sos_loop[0].somModel.cfg_dat_sel[1] = 1;
sos_loop[0].somModel.cfg_dat_vld[1] = 1;
sos_loop[0].somModel.cfg_miss_ptr[1] = 0;
sos_loop[0].somModel.tcam_data[2][0][0]=80'h00000000000000000000;
sos_loop[0].somModel.tcam_mask[2][0][0]=80'hffffffffffffffffffff;
sos_loop[0].somModel.tcam_data[2][1][0]=80'h00000000c76428a3ac18;
sos_loop[0].somModel.tcam_mask[2][1][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][2][0]=80'h000000006fa2b332a044;
sos_loop[0].somModel.tcam_mask[2][2][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][3][0]=80'h00000000df160ea7e244;
sos_loop[0].somModel.tcam_mask[2][3][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][4][0]=80'h00000000bde8a5158a2b;
sos_loop[0].somModel.tcam_mask[2][4][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][5][0]=80'h000000001c7fcaa5772f;
sos_loop[0].somModel.tcam_mask[2][5][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][6][0]=80'h00000000398bc2065413;
sos_loop[0].somModel.tcam_mask[2][6][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][7][0]=80'h00000000bf26a132d23e;
sos_loop[0].somModel.tcam_mask[2][7][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][8][0]=80'h000000002e5a52ddfb3f;
sos_loop[0].somModel.tcam_mask[2][8][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][9][0]=80'h000000000f9c4f448c4c;
sos_loop[0].somModel.tcam_mask[2][9][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][10][0]=80'h0000000035e4dd182f90;
sos_loop[0].somModel.tcam_mask[2][10][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][11][0]=80'h000000008513d0c50521;
sos_loop[0].somModel.tcam_mask[2][11][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][12][0]=80'h0000000035a66285b62e;
sos_loop[0].somModel.tcam_mask[2][12][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][13][0]=80'h000000004915d9de428f;
sos_loop[0].somModel.tcam_mask[2][13][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][14][0]=80'h000000003eff489073c2;
sos_loop[0].somModel.tcam_mask[2][14][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][15][0]=80'h00000000d00165db49c5;
sos_loop[0].somModel.tcam_mask[2][15][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][16][0]=80'h00000000c6e7d540048a;
sos_loop[0].somModel.tcam_mask[2][16][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][17][0]=80'h000000000d2cf31221e9;
sos_loop[0].somModel.tcam_mask[2][17][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][18][0]=80'h000000009cc2400c08bc;
sos_loop[0].somModel.tcam_mask[2][18][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][19][0]=80'h00000000e84ab68b1a24;
sos_loop[0].somModel.tcam_mask[2][19][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][20][0]=80'h00000000dc9c606e91ae;
sos_loop[0].somModel.tcam_mask[2][20][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][21][0]=80'h000000004b8ee53f7660;
sos_loop[0].somModel.tcam_mask[2][21][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][22][0]=80'h00000000a6dc109cdbbd;
sos_loop[0].somModel.tcam_mask[2][22][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][23][0]=80'h000000002e5acd726cb2;
sos_loop[0].somModel.tcam_mask[2][23][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][24][0]=80'h00000000bb30b2ecd487;
sos_loop[0].somModel.tcam_mask[2][24][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][25][0]=80'h000000009aeec82f8fac;
sos_loop[0].somModel.tcam_mask[2][25][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][26][0]=80'h00000000ab83fe2b985c;
sos_loop[0].somModel.tcam_mask[2][26][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][27][0]=80'h00000000ca3daac02b2f;
sos_loop[0].somModel.tcam_mask[2][27][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][28][0]=80'h000000001a893b2ffa10;
sos_loop[0].somModel.tcam_mask[2][28][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][29][0]=80'h00000000cb1ab883d9ca;
sos_loop[0].somModel.tcam_mask[2][29][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][30][0]=80'h000000006ddb0412e88d;
sos_loop[0].somModel.tcam_mask[2][30][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][31][0]=80'h0000000025d034a677c8;
sos_loop[0].somModel.tcam_mask[2][31][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][32][0]=80'h0000000002ee63ce89af;
sos_loop[0].somModel.tcam_mask[2][32][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[2][33][0]=80'h000000001ab5a710d843;
sos_loop[0].somModel.tcam_mask[2][33][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][34][0]=80'h0000000097e8c062f084;
sos_loop[0].somModel.tcam_mask[2][34][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][35][0]=80'h0000000030a809743d4f;
sos_loop[0].somModel.tcam_mask[2][35][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][36][0]=80'h0000000022420da7f8f4;
sos_loop[0].somModel.tcam_mask[2][36][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][37][0]=80'h00000000afaf284ad3bc;
sos_loop[0].somModel.tcam_mask[2][37][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][38][0]=80'h0000000053bd4f0d7794;
sos_loop[0].somModel.tcam_mask[2][38][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][39][0]=80'h000000005c0d39f2f061;
sos_loop[0].somModel.tcam_mask[2][39][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][40][0]=80'h000000009419a7ce074a;
sos_loop[0].somModel.tcam_mask[2][40][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][41][0]=80'h00000000052d45cc1e4a;
sos_loop[0].somModel.tcam_mask[2][41][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][42][0]=80'h000000009b30665b9971;
sos_loop[0].somModel.tcam_mask[2][42][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][43][0]=80'h0000000020d936f412c1;
sos_loop[0].somModel.tcam_mask[2][43][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][44][0]=80'h000000008b889af41550;
sos_loop[0].somModel.tcam_mask[2][44][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][45][0]=80'h00000000f91ce85e797d;
sos_loop[0].somModel.tcam_mask[2][45][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][46][0]=80'h0000000006e1dbd81191;
sos_loop[0].somModel.tcam_mask[2][46][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][47][0]=80'h00000000345e3c5f1365;
sos_loop[0].somModel.tcam_mask[2][47][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][48][0]=80'h000000008dceefe91dc9;
sos_loop[0].somModel.tcam_mask[2][48][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][49][0]=80'h00000000d47d2191ffed;
sos_loop[0].somModel.tcam_mask[2][49][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][50][0]=80'h000000007d341fbc821b;
sos_loop[0].somModel.tcam_mask[2][50][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][51][0]=80'h000000002e1c5d9ff7d9;
sos_loop[0].somModel.tcam_mask[2][51][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][52][0]=80'h00000000b7c667fd0324;
sos_loop[0].somModel.tcam_mask[2][52][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][53][0]=80'h000000004933bf21a16c;
sos_loop[0].somModel.tcam_mask[2][53][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][54][0]=80'h00000000f9724902347e;
sos_loop[0].somModel.tcam_mask[2][54][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][55][0]=80'h00000000aeb766b220db;
sos_loop[0].somModel.tcam_mask[2][55][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][56][0]=80'h00000000dbbc2a3224ab;
sos_loop[0].somModel.tcam_mask[2][56][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][57][0]=80'h00000000365a679e8085;
sos_loop[0].somModel.tcam_mask[2][57][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][58][0]=80'h00000000eeff7c2b7b33;
sos_loop[0].somModel.tcam_mask[2][58][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][59][0]=80'h0000000045bb6a31bb68;
sos_loop[0].somModel.tcam_mask[2][59][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][60][0]=80'h000000001a81b1c43f91;
sos_loop[0].somModel.tcam_mask[2][60][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][61][0]=80'h000000001de0ad29184a;
sos_loop[0].somModel.tcam_mask[2][61][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][62][0]=80'h000000004eb9229cd415;
sos_loop[0].somModel.tcam_mask[2][62][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][63][0]=80'h0000000075c39cfd15db;
sos_loop[0].somModel.tcam_mask[2][63][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][64][0]=80'h000000000bd7d9ddf726;
sos_loop[0].somModel.tcam_mask[2][64][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][65][0]=80'h00000000788ece7eed43;
sos_loop[0].somModel.tcam_mask[2][65][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][66][0]=80'h00000000689790000fff;
sos_loop[0].somModel.tcam_mask[2][66][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][67][0]=80'h0000000030fca31cf96b;
sos_loop[0].somModel.tcam_mask[2][67][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][68][0]=80'h00000000358975cc2823;
sos_loop[0].somModel.tcam_mask[2][68][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][69][0]=80'h000000006b1cd921c79d;
sos_loop[0].somModel.tcam_mask[2][69][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][70][0]=80'h00000000549a31ff63b7;
sos_loop[0].somModel.tcam_mask[2][70][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][71][0]=80'h00000000310dee607220;
sos_loop[0].somModel.tcam_mask[2][71][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][72][0]=80'h00000000af90fc2fb606;
sos_loop[0].somModel.tcam_mask[2][72][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][73][0]=80'h000000000db655000d3a;
sos_loop[0].somModel.tcam_mask[2][73][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][74][0]=80'h000000008bf35344ab45;
sos_loop[0].somModel.tcam_mask[2][74][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][75][0]=80'h000000002d8a38190b20;
sos_loop[0].somModel.tcam_mask[2][75][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][76][0]=80'h000000000263f7f66582;
sos_loop[0].somModel.tcam_mask[2][76][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[2][77][0]=80'h000000004dfc2ba4768d;
sos_loop[0].somModel.tcam_mask[2][77][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][78][0]=80'h00000000849983bfbe7a;
sos_loop[0].somModel.tcam_mask[2][78][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][79][0]=80'h000000001efcb2f4dd4d;
sos_loop[0].somModel.tcam_mask[2][79][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][80][0]=80'h0000000061e5a9de4569;
sos_loop[0].somModel.tcam_mask[2][80][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][81][0]=80'h00000000770c1c4bd3a5;
sos_loop[0].somModel.tcam_mask[2][81][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][82][0]=80'h00000000500562660aff;
sos_loop[0].somModel.tcam_mask[2][82][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][83][0]=80'h00000000a72a189143e2;
sos_loop[0].somModel.tcam_mask[2][83][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][84][0]=80'h0000000051a64abf0e09;
sos_loop[0].somModel.tcam_mask[2][84][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][85][0]=80'h000000001f5700abe928;
sos_loop[0].somModel.tcam_mask[2][85][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][86][0]=80'h00000000512e72fad6a2;
sos_loop[0].somModel.tcam_mask[2][86][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][87][0]=80'h000000005f3a530396cf;
sos_loop[0].somModel.tcam_mask[2][87][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][88][0]=80'h00000000748487400445;
sos_loop[0].somModel.tcam_mask[2][88][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][89][0]=80'h0000000087719fb3f864;
sos_loop[0].somModel.tcam_mask[2][89][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][90][0]=80'h00000000e88c8f60061d;
sos_loop[0].somModel.tcam_mask[2][90][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][91][0]=80'h000000009f6cc5f93019;
sos_loop[0].somModel.tcam_mask[2][91][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][92][0]=80'h00000000fa9df2c0fa11;
sos_loop[0].somModel.tcam_mask[2][92][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][93][0]=80'h000000003e5de237f4f3;
sos_loop[0].somModel.tcam_mask[2][93][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][94][0]=80'h000000001220e6f8b9fd;
sos_loop[0].somModel.tcam_mask[2][94][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][95][0]=80'h00000000ceb0c2f94c3c;
sos_loop[0].somModel.tcam_mask[2][95][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][96][0]=80'h000000001845b8356ded;
sos_loop[0].somModel.tcam_mask[2][96][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][97][0]=80'h00000000cb7d6f052ed9;
sos_loop[0].somModel.tcam_mask[2][97][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][98][0]=80'h00000000a1d827523dc7;
sos_loop[0].somModel.tcam_mask[2][98][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][99][0]=80'h000000000caf8264a3ea;
sos_loop[0].somModel.tcam_mask[2][99][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][100][0]=80'h0000000038ead3f12916;
sos_loop[0].somModel.tcam_mask[2][100][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][101][0]=80'h0000000013d2ee37c448;
sos_loop[0].somModel.tcam_mask[2][101][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][102][0]=80'h000000003c2fe7d9f34c;
sos_loop[0].somModel.tcam_mask[2][102][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][103][0]=80'h000000003c1db8626079;
sos_loop[0].somModel.tcam_mask[2][103][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][104][0]=80'h00000000865b861ca607;
sos_loop[0].somModel.tcam_mask[2][104][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][105][0]=80'h00000000794600c6d0f4;
sos_loop[0].somModel.tcam_mask[2][105][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][106][0]=80'h00000000e00c57f6e0b3;
sos_loop[0].somModel.tcam_mask[2][106][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][107][0]=80'h00000000e29db65e8903;
sos_loop[0].somModel.tcam_mask[2][107][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][108][0]=80'h000000008e261e6170f3;
sos_loop[0].somModel.tcam_mask[2][108][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][109][0]=80'h0000000066939b10ec73;
sos_loop[0].somModel.tcam_mask[2][109][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][110][0]=80'h0000000070c2e9c3c8eb;
sos_loop[0].somModel.tcam_mask[2][110][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][111][0]=80'h0000000045c66be84cf4;
sos_loop[0].somModel.tcam_mask[2][111][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][112][0]=80'h00000000232cef211d0e;
sos_loop[0].somModel.tcam_mask[2][112][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][113][0]=80'h0000000080542dda5aa2;
sos_loop[0].somModel.tcam_mask[2][113][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][114][0]=80'h00000000474effbc30dd;
sos_loop[0].somModel.tcam_mask[2][114][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][115][0]=80'h00000000e4cebd5c6fa4;
sos_loop[0].somModel.tcam_mask[2][115][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][116][0]=80'h00000000af6a54830375;
sos_loop[0].somModel.tcam_mask[2][116][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][117][0]=80'h000000008ef028be44c1;
sos_loop[0].somModel.tcam_mask[2][117][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][118][0]=80'h000000005fdca8436bf4;
sos_loop[0].somModel.tcam_mask[2][118][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][119][0]=80'h000000006e7e1c15bd08;
sos_loop[0].somModel.tcam_mask[2][119][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][120][0]=80'h00000000134c1f65fd66;
sos_loop[0].somModel.tcam_mask[2][120][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][121][0]=80'h00000000cea87493679f;
sos_loop[0].somModel.tcam_mask[2][121][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][122][0]=80'h00000000ceb7bc309c1a;
sos_loop[0].somModel.tcam_mask[2][122][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][123][0]=80'h0000000061a6f8771878;
sos_loop[0].somModel.tcam_mask[2][123][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][124][0]=80'h00000000cedef6a567fe;
sos_loop[0].somModel.tcam_mask[2][124][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][125][0]=80'h000000002e32a08622cd;
sos_loop[0].somModel.tcam_mask[2][125][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][126][0]=80'h000000005356e16b8fd7;
sos_loop[0].somModel.tcam_mask[2][126][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][127][0]=80'h00000000fd605bd942c3;
sos_loop[0].somModel.tcam_mask[2][127][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][128][0]=80'h0000000000d5f103f449;
sos_loop[0].somModel.tcam_mask[2][128][0]=80'hffffffffff0000000000;
sos_loop[0].somModel.tcam_data[2][129][0]=80'h000000005f57f4362b22;
sos_loop[0].somModel.tcam_mask[2][129][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][130][0]=80'h000000002e67f284f871;
sos_loop[0].somModel.tcam_mask[2][130][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][131][0]=80'h00000000ecd79dcadc01;
sos_loop[0].somModel.tcam_mask[2][131][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][132][0]=80'h00000000e00525c7b0f8;
sos_loop[0].somModel.tcam_mask[2][132][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][133][0]=80'h00000000b3cf483e6c80;
sos_loop[0].somModel.tcam_mask[2][133][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][134][0]=80'h0000000077eb26f31bbe;
sos_loop[0].somModel.tcam_mask[2][134][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][135][0]=80'h000000008b676c49d915;
sos_loop[0].somModel.tcam_mask[2][135][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][136][0]=80'h000000000a2822acbd35;
sos_loop[0].somModel.tcam_mask[2][136][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][137][0]=80'h0000000003a257929df1;
sos_loop[0].somModel.tcam_mask[2][137][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[2][138][0]=80'h00000000e9b0e1c40a18;
sos_loop[0].somModel.tcam_mask[2][138][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][139][0]=80'h000000003f10a0b32f42;
sos_loop[0].somModel.tcam_mask[2][139][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][140][0]=80'h00000000f8a042a8b1d1;
sos_loop[0].somModel.tcam_mask[2][140][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][141][0]=80'h00000000c010041f98fe;
sos_loop[0].somModel.tcam_mask[2][141][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][142][0]=80'h000000006f5155d6bf2a;
sos_loop[0].somModel.tcam_mask[2][142][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][143][0]=80'h000000006174e0aee88e;
sos_loop[0].somModel.tcam_mask[2][143][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][144][0]=80'h00000000d8f296505931;
sos_loop[0].somModel.tcam_mask[2][144][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][145][0]=80'h00000000e512e3c64789;
sos_loop[0].somModel.tcam_mask[2][145][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][146][0]=80'h00000000373e0b9976b9;
sos_loop[0].somModel.tcam_mask[2][146][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][147][0]=80'h0000000003e7dacda18b;
sos_loop[0].somModel.tcam_mask[2][147][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[2][148][0]=80'h000000000964ddbc00a5;
sos_loop[0].somModel.tcam_mask[2][148][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][149][0]=80'h0000000054781b947c65;
sos_loop[0].somModel.tcam_mask[2][149][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][150][0]=80'h000000004e476ae23070;
sos_loop[0].somModel.tcam_mask[2][150][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][151][0]=80'h00000000965a202c5dd1;
sos_loop[0].somModel.tcam_mask[2][151][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][152][0]=80'h000000006eeef25e5a0e;
sos_loop[0].somModel.tcam_mask[2][152][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][153][0]=80'h00000000bd9be825e53c;
sos_loop[0].somModel.tcam_mask[2][153][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][154][0]=80'h000000005a0d2b0e2652;
sos_loop[0].somModel.tcam_mask[2][154][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][155][0]=80'h00000000f02c2960a78f;
sos_loop[0].somModel.tcam_mask[2][155][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][156][0]=80'h0000000043801573ed5c;
sos_loop[0].somModel.tcam_mask[2][156][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][157][0]=80'h0000000034d1a3628645;
sos_loop[0].somModel.tcam_mask[2][157][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][158][0]=80'h00000000476d2c7ebc16;
sos_loop[0].somModel.tcam_mask[2][158][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][159][0]=80'h00000000a17de6c9b9c6;
sos_loop[0].somModel.tcam_mask[2][159][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][160][0]=80'h000000002e3b2da7cb0e;
sos_loop[0].somModel.tcam_mask[2][160][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][161][0]=80'h00000000618fe75b3a00;
sos_loop[0].somModel.tcam_mask[2][161][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][162][0]=80'h000000007868e9b929a2;
sos_loop[0].somModel.tcam_mask[2][162][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][163][0]=80'h00000000cbe5e4137d1a;
sos_loop[0].somModel.tcam_mask[2][163][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][164][0]=80'h000000006771e8c490b5;
sos_loop[0].somModel.tcam_mask[2][164][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][165][0]=80'h000000007be9cc15dbad;
sos_loop[0].somModel.tcam_mask[2][165][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][166][0]=80'h000000008c89b097b14c;
sos_loop[0].somModel.tcam_mask[2][166][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][167][0]=80'h00000000f2124342ae18;
sos_loop[0].somModel.tcam_mask[2][167][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][168][0]=80'h00000000330261ba3670;
sos_loop[0].somModel.tcam_mask[2][168][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][169][0]=80'h0000000042c4edb6d896;
sos_loop[0].somModel.tcam_mask[2][169][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][170][0]=80'h0000000023a570bc32da;
sos_loop[0].somModel.tcam_mask[2][170][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][171][0]=80'h00000000db4f2973fc73;
sos_loop[0].somModel.tcam_mask[2][171][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][172][0]=80'h000000004c40d88318b1;
sos_loop[0].somModel.tcam_mask[2][172][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][173][0]=80'h000000001273739101e3;
sos_loop[0].somModel.tcam_mask[2][173][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][174][0]=80'h000000009c2ebac8770d;
sos_loop[0].somModel.tcam_mask[2][174][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][175][0]=80'h00000000aaeaffde1744;
sos_loop[0].somModel.tcam_mask[2][175][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][176][0]=80'h0000000067b1d0406ac4;
sos_loop[0].somModel.tcam_mask[2][176][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][177][0]=80'h00000000602be7c25423;
sos_loop[0].somModel.tcam_mask[2][177][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][178][0]=80'h000000007bd2374d89da;
sos_loop[0].somModel.tcam_mask[2][178][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][179][0]=80'h00000000484efbf68ee5;
sos_loop[0].somModel.tcam_mask[2][179][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][180][0]=80'h000000008c2970d5df55;
sos_loop[0].somModel.tcam_mask[2][180][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][181][0]=80'h00000000aec65cebfe7b;
sos_loop[0].somModel.tcam_mask[2][181][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][182][0]=80'h0000000094dfc4cad63a;
sos_loop[0].somModel.tcam_mask[2][182][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][183][0]=80'h0000000016398c9c5329;
sos_loop[0].somModel.tcam_mask[2][183][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][184][0]=80'h00000000c1d9c5b84501;
sos_loop[0].somModel.tcam_mask[2][184][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][185][0]=80'h00000000d1ad3332662b;
sos_loop[0].somModel.tcam_mask[2][185][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][186][0]=80'h00000000b91d094ca5fa;
sos_loop[0].somModel.tcam_mask[2][186][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][187][0]=80'h0000000066807169ce5b;
sos_loop[0].somModel.tcam_mask[2][187][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][188][0]=80'h000000006ef096e4f564;
sos_loop[0].somModel.tcam_mask[2][188][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][189][0]=80'h00000000328864e675f7;
sos_loop[0].somModel.tcam_mask[2][189][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][190][0]=80'h000000007dae2b0e1b45;
sos_loop[0].somModel.tcam_mask[2][190][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][191][0]=80'h00000000bcb94b47b6e1;
sos_loop[0].somModel.tcam_mask[2][191][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][192][0]=80'h00000000969630df4be5;
sos_loop[0].somModel.tcam_mask[2][192][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][193][0]=80'h000000008fa1021a531a;
sos_loop[0].somModel.tcam_mask[2][193][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][194][0]=80'h00000000872d61d5debf;
sos_loop[0].somModel.tcam_mask[2][194][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][195][0]=80'h00000000991610788933;
sos_loop[0].somModel.tcam_mask[2][195][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][196][0]=80'h000000000abf899e0a35;
sos_loop[0].somModel.tcam_mask[2][196][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][197][0]=80'h000000009a50b37b4c4e;
sos_loop[0].somModel.tcam_mask[2][197][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][198][0]=80'h00000000a57859f9c477;
sos_loop[0].somModel.tcam_mask[2][198][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][199][0]=80'h000000000079cd60c49c;
sos_loop[0].somModel.tcam_mask[2][199][0]=80'hffffffffff8000000000;
sos_loop[0].somModel.tcam_data[2][200][0]=80'h00000000116a5a1abd7d;
sos_loop[0].somModel.tcam_mask[2][200][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][201][0]=80'h00000000c21fd0b46818;
sos_loop[0].somModel.tcam_mask[2][201][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][202][0]=80'h00000000cb7c1d8cfffa;
sos_loop[0].somModel.tcam_mask[2][202][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][203][0]=80'h000000005da2668e789f;
sos_loop[0].somModel.tcam_mask[2][203][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][204][0]=80'h00000000a975554d1660;
sos_loop[0].somModel.tcam_mask[2][204][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][205][0]=80'h00000000f527f8412a24;
sos_loop[0].somModel.tcam_mask[2][205][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][206][0]=80'h000000006e7cabe12a47;
sos_loop[0].somModel.tcam_mask[2][206][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][207][0]=80'h00000000ecce1c4cd86e;
sos_loop[0].somModel.tcam_mask[2][207][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][208][0]=80'h0000000072d3d3fcd72b;
sos_loop[0].somModel.tcam_mask[2][208][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][209][0]=80'h00000000839e1fb55d44;
sos_loop[0].somModel.tcam_mask[2][209][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][210][0]=80'h00000000478398e0b9ee;
sos_loop[0].somModel.tcam_mask[2][210][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][211][0]=80'h000000008530d50e759f;
sos_loop[0].somModel.tcam_mask[2][211][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][212][0]=80'h0000000011f968361ebd;
sos_loop[0].somModel.tcam_mask[2][212][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][213][0]=80'h000000008ce994cc083f;
sos_loop[0].somModel.tcam_mask[2][213][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][214][0]=80'h000000002c23f84988ee;
sos_loop[0].somModel.tcam_mask[2][214][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][215][0]=80'h000000009760938f25c2;
sos_loop[0].somModel.tcam_mask[2][215][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][216][0]=80'h00000000274efbfa8211;
sos_loop[0].somModel.tcam_mask[2][216][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][217][0]=80'h00000000694132b93ba3;
sos_loop[0].somModel.tcam_mask[2][217][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][218][0]=80'h000000000682f3056401;
sos_loop[0].somModel.tcam_mask[2][218][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][219][0]=80'h00000000d1c36a785d4f;
sos_loop[0].somModel.tcam_mask[2][219][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][220][0]=80'h000000004ae9b6d2ef4f;
sos_loop[0].somModel.tcam_mask[2][220][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][221][0]=80'h00000000c9c32ab41eeb;
sos_loop[0].somModel.tcam_mask[2][221][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][222][0]=80'h00000000cbc076ebe28e;
sos_loop[0].somModel.tcam_mask[2][222][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][223][0]=80'h00000000fbda31fd76c0;
sos_loop[0].somModel.tcam_mask[2][223][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][224][0]=80'h000000009a099a151b35;
sos_loop[0].somModel.tcam_mask[2][224][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][225][0]=80'h0000000054a1681b3ffb;
sos_loop[0].somModel.tcam_mask[2][225][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][226][0]=80'h00000000f0cf8f9ee272;
sos_loop[0].somModel.tcam_mask[2][226][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][227][0]=80'h000000003f535b44d28a;
sos_loop[0].somModel.tcam_mask[2][227][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][228][0]=80'h000000007ae44fa333c8;
sos_loop[0].somModel.tcam_mask[2][228][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][229][0]=80'h00000000b665ce7f735a;
sos_loop[0].somModel.tcam_mask[2][229][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][230][0]=80'h00000000626c7ae8774d;
sos_loop[0].somModel.tcam_mask[2][230][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][231][0]=80'h00000000f3cddb51d392;
sos_loop[0].somModel.tcam_mask[2][231][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][232][0]=80'h00000000944a75a8319c;
sos_loop[0].somModel.tcam_mask[2][232][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][233][0]=80'h00000000eaacb9890fae;
sos_loop[0].somModel.tcam_mask[2][233][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][234][0]=80'h00000000046f6540ec7f;
sos_loop[0].somModel.tcam_mask[2][234][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][235][0]=80'h00000000c6088fc1bd3d;
sos_loop[0].somModel.tcam_mask[2][235][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][236][0]=80'h000000005e0b61c56031;
sos_loop[0].somModel.tcam_mask[2][236][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][237][0]=80'h00000000027b4c51c3bb;
sos_loop[0].somModel.tcam_mask[2][237][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[2][238][0]=80'h00000000be4d82d7e60e;
sos_loop[0].somModel.tcam_mask[2][238][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][239][0]=80'h000000007eef6a0932c5;
sos_loop[0].somModel.tcam_mask[2][239][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][240][0]=80'h00000000564f40cb3bc6;
sos_loop[0].somModel.tcam_mask[2][240][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][241][0]=80'h0000000049ba0e14ede1;
sos_loop[0].somModel.tcam_mask[2][241][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][242][0]=80'h000000000ffa1385e8e1;
sos_loop[0].somModel.tcam_mask[2][242][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][243][0]=80'h00000000c2a6a6c5875c;
sos_loop[0].somModel.tcam_mask[2][243][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][244][0]=80'h0000000046ed88992ff9;
sos_loop[0].somModel.tcam_mask[2][244][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][245][0]=80'h000000007bd52c488741;
sos_loop[0].somModel.tcam_mask[2][245][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][246][0]=80'h00000000dd037b320186;
sos_loop[0].somModel.tcam_mask[2][246][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][247][0]=80'h00000000bc45bae8ac0a;
sos_loop[0].somModel.tcam_mask[2][247][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][248][0]=80'h000000005b06c7e96f30;
sos_loop[0].somModel.tcam_mask[2][248][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][249][0]=80'h00000000d4ddc557a673;
sos_loop[0].somModel.tcam_mask[2][249][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][250][0]=80'h0000000053ec21af6aa7;
sos_loop[0].somModel.tcam_mask[2][250][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][251][0]=80'h0000000017ac57f88e87;
sos_loop[0].somModel.tcam_mask[2][251][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][252][0]=80'h00000000a4100e4032cc;
sos_loop[0].somModel.tcam_mask[2][252][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][253][0]=80'h00000000140fa51dda60;
sos_loop[0].somModel.tcam_mask[2][253][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][254][0]=80'h00000000ba76b63b04af;
sos_loop[0].somModel.tcam_mask[2][254][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][255][0]=80'h000000007bf30212d42d;
sos_loop[0].somModel.tcam_mask[2][255][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][256][0]=80'h00000000389a856d0929;
sos_loop[0].somModel.tcam_mask[2][256][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][257][0]=80'h00000000971def77bfa0;
sos_loop[0].somModel.tcam_mask[2][257][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][258][0]=80'h000000007fea6ca2dda9;
sos_loop[0].somModel.tcam_mask[2][258][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][259][0]=80'h000000006cc87b7163e1;
sos_loop[0].somModel.tcam_mask[2][259][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][260][0]=80'h00000000652f37432033;
sos_loop[0].somModel.tcam_mask[2][260][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][261][0]=80'h0000000094ca0afeaf40;
sos_loop[0].somModel.tcam_mask[2][261][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][262][0]=80'h00000000aa6075a82cfd;
sos_loop[0].somModel.tcam_mask[2][262][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][263][0]=80'h00000000e393132fbd4d;
sos_loop[0].somModel.tcam_mask[2][263][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][264][0]=80'h000000008617fb8769a3;
sos_loop[0].somModel.tcam_mask[2][264][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][265][0]=80'h00000000d45704f554fa;
sos_loop[0].somModel.tcam_mask[2][265][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][266][0]=80'h00000000083aeac67707;
sos_loop[0].somModel.tcam_mask[2][266][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][267][0]=80'h00000000ad11dd592c9a;
sos_loop[0].somModel.tcam_mask[2][267][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][268][0]=80'h00000000199fcd09ed28;
sos_loop[0].somModel.tcam_mask[2][268][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][269][0]=80'h00000000306fc67d4fd2;
sos_loop[0].somModel.tcam_mask[2][269][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][270][0]=80'h00000000ded308236673;
sos_loop[0].somModel.tcam_mask[2][270][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][271][0]=80'h000000006bb4f3981543;
sos_loop[0].somModel.tcam_mask[2][271][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][272][0]=80'h0000000028d774fa8bab;
sos_loop[0].somModel.tcam_mask[2][272][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][273][0]=80'h000000005f39e126fa40;
sos_loop[0].somModel.tcam_mask[2][273][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][274][0]=80'h000000004ec1930dd830;
sos_loop[0].somModel.tcam_mask[2][274][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][275][0]=80'h000000002eabafa47444;
sos_loop[0].somModel.tcam_mask[2][275][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][276][0]=80'h00000000f2c4354979b5;
sos_loop[0].somModel.tcam_mask[2][276][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][277][0]=80'h000000004375ff2839ff;
sos_loop[0].somModel.tcam_mask[2][277][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][278][0]=80'h00000000831847d750e3;
sos_loop[0].somModel.tcam_mask[2][278][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][279][0]=80'h000000006d4ff70a7fc3;
sos_loop[0].somModel.tcam_mask[2][279][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][280][0]=80'h0000000067633ad96690;
sos_loop[0].somModel.tcam_mask[2][280][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][281][0]=80'h0000000058b1bb7ab35b;
sos_loop[0].somModel.tcam_mask[2][281][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][282][0]=80'h00000000378d65b1297a;
sos_loop[0].somModel.tcam_mask[2][282][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][283][0]=80'h000000008ab24a720a34;
sos_loop[0].somModel.tcam_mask[2][283][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][284][0]=80'h000000009b617faf808a;
sos_loop[0].somModel.tcam_mask[2][284][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][285][0]=80'h000000002b5be33345f9;
sos_loop[0].somModel.tcam_mask[2][285][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][286][0]=80'h0000000080b069925240;
sos_loop[0].somModel.tcam_mask[2][286][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][287][0]=80'h0000000064819ae5ce38;
sos_loop[0].somModel.tcam_mask[2][287][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][288][0]=80'h00000000c8a2886319ad;
sos_loop[0].somModel.tcam_mask[2][288][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][289][0]=80'h00000000bba80680cd74;
sos_loop[0].somModel.tcam_mask[2][289][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][290][0]=80'h00000000c624c1780420;
sos_loop[0].somModel.tcam_mask[2][290][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][291][0]=80'h000000000df4dc19f8a0;
sos_loop[0].somModel.tcam_mask[2][291][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][292][0]=80'h00000000bf4fc4c5109d;
sos_loop[0].somModel.tcam_mask[2][292][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][293][0]=80'h00000000230e53a6e40d;
sos_loop[0].somModel.tcam_mask[2][293][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][294][0]=80'h000000006a8845704812;
sos_loop[0].somModel.tcam_mask[2][294][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][295][0]=80'h00000000d02d7e61c3ff;
sos_loop[0].somModel.tcam_mask[2][295][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][296][0]=80'h0000000042d9ad4b7cb5;
sos_loop[0].somModel.tcam_mask[2][296][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][297][0]=80'h000000006620c43e40cd;
sos_loop[0].somModel.tcam_mask[2][297][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][298][0]=80'h00000000572b2a5075a9;
sos_loop[0].somModel.tcam_mask[2][298][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][299][0]=80'h000000000bc0a3cd8632;
sos_loop[0].somModel.tcam_mask[2][299][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][300][0]=80'h00000000318840f45c23;
sos_loop[0].somModel.tcam_mask[2][300][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][301][0]=80'h000000007ec0b9f2df84;
sos_loop[0].somModel.tcam_mask[2][301][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][302][0]=80'h000000000708eaeea371;
sos_loop[0].somModel.tcam_mask[2][302][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][303][0]=80'h0000000029e3e9901c1f;
sos_loop[0].somModel.tcam_mask[2][303][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][304][0]=80'h00000000f4f0fb40376f;
sos_loop[0].somModel.tcam_mask[2][304][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][305][0]=80'h000000007de8c27c7bf8;
sos_loop[0].somModel.tcam_mask[2][305][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][306][0]=80'h00000000722214538bb3;
sos_loop[0].somModel.tcam_mask[2][306][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][307][0]=80'h00000000b35284a2e8f3;
sos_loop[0].somModel.tcam_mask[2][307][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][308][0]=80'h00000000c1e963dc4088;
sos_loop[0].somModel.tcam_mask[2][308][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][309][0]=80'h0000000050d5503770e6;
sos_loop[0].somModel.tcam_mask[2][309][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][310][0]=80'h00000000b63951662a30;
sos_loop[0].somModel.tcam_mask[2][310][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][311][0]=80'h000000007eddea567619;
sos_loop[0].somModel.tcam_mask[2][311][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][312][0]=80'h000000004eab0a109e8f;
sos_loop[0].somModel.tcam_mask[2][312][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][313][0]=80'h00000000e549f26a551a;
sos_loop[0].somModel.tcam_mask[2][313][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][314][0]=80'h00000000161e12d7d5f4;
sos_loop[0].somModel.tcam_mask[2][314][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][315][0]=80'h000000002fb8691cf03d;
sos_loop[0].somModel.tcam_mask[2][315][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][316][0]=80'h000000006d0dd414bd88;
sos_loop[0].somModel.tcam_mask[2][316][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][317][0]=80'h00000000d47f0cfd8269;
sos_loop[0].somModel.tcam_mask[2][317][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][318][0]=80'h00000000e7fe58f76aac;
sos_loop[0].somModel.tcam_mask[2][318][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][319][0]=80'h00000000cddb5437e4b9;
sos_loop[0].somModel.tcam_mask[2][319][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][320][0]=80'h0000000058ac2d7d65c1;
sos_loop[0].somModel.tcam_mask[2][320][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][321][0]=80'h00000000e81d8eb85034;
sos_loop[0].somModel.tcam_mask[2][321][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][322][0]=80'h00000000a6fb99d69d1b;
sos_loop[0].somModel.tcam_mask[2][322][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][323][0]=80'h0000000085db0f2ad52e;
sos_loop[0].somModel.tcam_mask[2][323][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][324][0]=80'h00000000ba447f49c0b1;
sos_loop[0].somModel.tcam_mask[2][324][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][325][0]=80'h0000000099d3496acd35;
sos_loop[0].somModel.tcam_mask[2][325][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][326][0]=80'h0000000040e7e1b07303;
sos_loop[0].somModel.tcam_mask[2][326][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][327][0]=80'h0000000055f948ebe91d;
sos_loop[0].somModel.tcam_mask[2][327][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][328][0]=80'h00000000392c0459ce02;
sos_loop[0].somModel.tcam_mask[2][328][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][329][0]=80'h000000007e3d419f5d34;
sos_loop[0].somModel.tcam_mask[2][329][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][330][0]=80'h00000000e74efb58eaa7;
sos_loop[0].somModel.tcam_mask[2][330][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][331][0]=80'h00000000f83f581e4482;
sos_loop[0].somModel.tcam_mask[2][331][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][332][0]=80'h000000009cce1dfeef14;
sos_loop[0].somModel.tcam_mask[2][332][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][333][0]=80'h000000004b70936e9f64;
sos_loop[0].somModel.tcam_mask[2][333][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][334][0]=80'h000000008f60bf446783;
sos_loop[0].somModel.tcam_mask[2][334][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][335][0]=80'h0000000093a9046448e2;
sos_loop[0].somModel.tcam_mask[2][335][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][336][0]=80'h000000006e3ce4ac6730;
sos_loop[0].somModel.tcam_mask[2][336][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][337][0]=80'h0000000084de22fbc40a;
sos_loop[0].somModel.tcam_mask[2][337][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][338][0]=80'h000000002d98732c0914;
sos_loop[0].somModel.tcam_mask[2][338][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][339][0]=80'h00000000588e0584287c;
sos_loop[0].somModel.tcam_mask[2][339][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][340][0]=80'h000000008f50e0497e89;
sos_loop[0].somModel.tcam_mask[2][340][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][341][0]=80'h00000000b0e119fb2555;
sos_loop[0].somModel.tcam_mask[2][341][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][342][0]=80'h000000004cd3c2cde21a;
sos_loop[0].somModel.tcam_mask[2][342][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][343][0]=80'h00000000da342cb3beee;
sos_loop[0].somModel.tcam_mask[2][343][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][344][0]=80'h000000009f7fc5e6a042;
sos_loop[0].somModel.tcam_mask[2][344][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][345][0]=80'h00000000cc5300c82669;
sos_loop[0].somModel.tcam_mask[2][345][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][346][0]=80'h000000006a1ec386bf00;
sos_loop[0].somModel.tcam_mask[2][346][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][347][0]=80'h000000002317e8d90545;
sos_loop[0].somModel.tcam_mask[2][347][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][348][0]=80'h000000008d4fe98625cf;
sos_loop[0].somModel.tcam_mask[2][348][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][349][0]=80'h00000000060665e2c19e;
sos_loop[0].somModel.tcam_mask[2][349][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][350][0]=80'h00000000596674fbbfb1;
sos_loop[0].somModel.tcam_mask[2][350][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][351][0]=80'h000000005c7688d8aad5;
sos_loop[0].somModel.tcam_mask[2][351][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][352][0]=80'h0000000099c3cb202d30;
sos_loop[0].somModel.tcam_mask[2][352][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][353][0]=80'h00000000a86ac83a7681;
sos_loop[0].somModel.tcam_mask[2][353][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][354][0]=80'h00000000f9f330aaf7e5;
sos_loop[0].somModel.tcam_mask[2][354][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][355][0]=80'h000000003c3dcdb988e5;
sos_loop[0].somModel.tcam_mask[2][355][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][356][0]=80'h0000000082440e73e0a4;
sos_loop[0].somModel.tcam_mask[2][356][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][357][0]=80'h00000000deb63d376bdd;
sos_loop[0].somModel.tcam_mask[2][357][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][358][0]=80'h000000003f13c6d986da;
sos_loop[0].somModel.tcam_mask[2][358][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][359][0]=80'h00000000959a11161a8a;
sos_loop[0].somModel.tcam_mask[2][359][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][360][0]=80'h0000000004fc4b9709a2;
sos_loop[0].somModel.tcam_mask[2][360][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][361][0]=80'h000000000603260a4fa8;
sos_loop[0].somModel.tcam_mask[2][361][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][362][0]=80'h00000000317642426d30;
sos_loop[0].somModel.tcam_mask[2][362][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][363][0]=80'h0000000093eea5159da0;
sos_loop[0].somModel.tcam_mask[2][363][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][364][0]=80'h00000000a6a6c5effbb8;
sos_loop[0].somModel.tcam_mask[2][364][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][365][0]=80'h000000009a556fc0f1e1;
sos_loop[0].somModel.tcam_mask[2][365][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][366][0]=80'h00000000ca8bfde422b1;
sos_loop[0].somModel.tcam_mask[2][366][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][367][0]=80'h000000006b3d4da4a0e4;
sos_loop[0].somModel.tcam_mask[2][367][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][368][0]=80'h00000000b8725432eee0;
sos_loop[0].somModel.tcam_mask[2][368][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][369][0]=80'h000000002a5f4d97572c;
sos_loop[0].somModel.tcam_mask[2][369][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][370][0]=80'h0000000003f4b2f37c91;
sos_loop[0].somModel.tcam_mask[2][370][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[2][371][0]=80'h000000006d012a56f306;
sos_loop[0].somModel.tcam_mask[2][371][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][372][0]=80'h00000000f39c18ff7423;
sos_loop[0].somModel.tcam_mask[2][372][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][373][0]=80'h0000000064fe54c3d020;
sos_loop[0].somModel.tcam_mask[2][373][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][374][0]=80'h000000005941386df853;
sos_loop[0].somModel.tcam_mask[2][374][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][375][0]=80'h00000000fd5081a7023d;
sos_loop[0].somModel.tcam_mask[2][375][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][376][0]=80'h0000000059d252677e44;
sos_loop[0].somModel.tcam_mask[2][376][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][377][0]=80'h00000000b1ef710456c8;
sos_loop[0].somModel.tcam_mask[2][377][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][378][0]=80'h000000008a3b29afa55f;
sos_loop[0].somModel.tcam_mask[2][378][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][379][0]=80'h00000000a8f4af7c920a;
sos_loop[0].somModel.tcam_mask[2][379][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][380][0]=80'h000000009b5b556528f0;
sos_loop[0].somModel.tcam_mask[2][380][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][381][0]=80'h000000008d75c4ce6384;
sos_loop[0].somModel.tcam_mask[2][381][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][382][0]=80'h00000000644e172a4d39;
sos_loop[0].somModel.tcam_mask[2][382][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][383][0]=80'h000000004e2c31c4e9bf;
sos_loop[0].somModel.tcam_mask[2][383][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][384][0]=80'h00000000fb16e104670e;
sos_loop[0].somModel.tcam_mask[2][384][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][385][0]=80'h00000000edda66338267;
sos_loop[0].somModel.tcam_mask[2][385][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][386][0]=80'h00000000028c12a16f1b;
sos_loop[0].somModel.tcam_mask[2][386][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[2][387][0]=80'h00000000ff84824ad314;
sos_loop[0].somModel.tcam_mask[2][387][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][388][0]=80'h000000000be7756aeeab;
sos_loop[0].somModel.tcam_mask[2][388][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][389][0]=80'h000000007e61e055303f;
sos_loop[0].somModel.tcam_mask[2][389][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][390][0]=80'h00000000aac7193a22af;
sos_loop[0].somModel.tcam_mask[2][390][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][391][0]=80'h00000000565f0106873e;
sos_loop[0].somModel.tcam_mask[2][391][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][392][0]=80'h0000000075032e61802d;
sos_loop[0].somModel.tcam_mask[2][392][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][393][0]=80'h00000000f2f7c9dbbf6e;
sos_loop[0].somModel.tcam_mask[2][393][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][394][0]=80'h00000000c616b82074dc;
sos_loop[0].somModel.tcam_mask[2][394][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][395][0]=80'h000000009b90c73a26b9;
sos_loop[0].somModel.tcam_mask[2][395][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][396][0]=80'h00000000f1aad48501e0;
sos_loop[0].somModel.tcam_mask[2][396][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][397][0]=80'h00000000b50e5a5b2331;
sos_loop[0].somModel.tcam_mask[2][397][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][398][0]=80'h000000000536e70ff511;
sos_loop[0].somModel.tcam_mask[2][398][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][399][0]=80'h00000000500f137223d6;
sos_loop[0].somModel.tcam_mask[2][399][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][400][0]=80'h000000002791051b62a6;
sos_loop[0].somModel.tcam_mask[2][400][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][401][0]=80'h00000000c4eb2c045df0;
sos_loop[0].somModel.tcam_mask[2][401][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][402][0]=80'h00000000a4ad1b4e4c65;
sos_loop[0].somModel.tcam_mask[2][402][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][403][0]=80'h000000005dcd203c62ab;
sos_loop[0].somModel.tcam_mask[2][403][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][404][0]=80'h00000000bd2053fe1aa1;
sos_loop[0].somModel.tcam_mask[2][404][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][405][0]=80'h00000000dd873733eebd;
sos_loop[0].somModel.tcam_mask[2][405][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][406][0]=80'h00000000d5cc8944cc44;
sos_loop[0].somModel.tcam_mask[2][406][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][407][0]=80'h00000000df75e34c1d60;
sos_loop[0].somModel.tcam_mask[2][407][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][408][0]=80'h0000000069516c90e02b;
sos_loop[0].somModel.tcam_mask[2][408][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][409][0]=80'h00000000ba7434218648;
sos_loop[0].somModel.tcam_mask[2][409][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][410][0]=80'h0000000075995e082cc9;
sos_loop[0].somModel.tcam_mask[2][410][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][411][0]=80'h000000008f8a0618c492;
sos_loop[0].somModel.tcam_mask[2][411][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][412][0]=80'h0000000085652adefb50;
sos_loop[0].somModel.tcam_mask[2][412][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][413][0]=80'h0000000084e3bbb346a9;
sos_loop[0].somModel.tcam_mask[2][413][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][414][0]=80'h00000000ce288545ff5c;
sos_loop[0].somModel.tcam_mask[2][414][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][415][0]=80'h00000000f34840529bc7;
sos_loop[0].somModel.tcam_mask[2][415][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][416][0]=80'h0000000093b680734ca8;
sos_loop[0].somModel.tcam_mask[2][416][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][417][0]=80'h000000006d3e5930bf31;
sos_loop[0].somModel.tcam_mask[2][417][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][418][0]=80'h000000004c6bb4e13dd2;
sos_loop[0].somModel.tcam_mask[2][418][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][419][0]=80'h00000000c17e7cae146d;
sos_loop[0].somModel.tcam_mask[2][419][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][420][0]=80'h000000003a01e234f448;
sos_loop[0].somModel.tcam_mask[2][420][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][421][0]=80'h000000001f6089a70d31;
sos_loop[0].somModel.tcam_mask[2][421][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][422][0]=80'h00000000e9910acedf01;
sos_loop[0].somModel.tcam_mask[2][422][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][423][0]=80'h0000000092c1be63a45c;
sos_loop[0].somModel.tcam_mask[2][423][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][424][0]=80'h0000000077250b5545e8;
sos_loop[0].somModel.tcam_mask[2][424][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][425][0]=80'h0000000041875a4af1b4;
sos_loop[0].somModel.tcam_mask[2][425][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][426][0]=80'h000000001f7188b8f195;
sos_loop[0].somModel.tcam_mask[2][426][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][427][0]=80'h00000000e7043697f5e9;
sos_loop[0].somModel.tcam_mask[2][427][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][428][0]=80'h00000000ccb0a5325cbe;
sos_loop[0].somModel.tcam_mask[2][428][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][429][0]=80'h00000000f77c99d0ae10;
sos_loop[0].somModel.tcam_mask[2][429][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][430][0]=80'h0000000051c66267cec7;
sos_loop[0].somModel.tcam_mask[2][430][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][431][0]=80'h00000000a3eb7b517f7d;
sos_loop[0].somModel.tcam_mask[2][431][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][432][0]=80'h000000005e4b84a9a324;
sos_loop[0].somModel.tcam_mask[2][432][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][433][0]=80'h00000000263366d9a934;
sos_loop[0].somModel.tcam_mask[2][433][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][434][0]=80'h0000000035cd167e2bad;
sos_loop[0].somModel.tcam_mask[2][434][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][435][0]=80'h000000000b2c3bbf8fba;
sos_loop[0].somModel.tcam_mask[2][435][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][436][0]=80'h000000008f19a66976c7;
sos_loop[0].somModel.tcam_mask[2][436][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][437][0]=80'h00000000e0b42c35622b;
sos_loop[0].somModel.tcam_mask[2][437][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][438][0]=80'h00000000dca9a6f1782c;
sos_loop[0].somModel.tcam_mask[2][438][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][439][0]=80'h000000009a1541c274a2;
sos_loop[0].somModel.tcam_mask[2][439][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][440][0]=80'h0000000044768a38b95d;
sos_loop[0].somModel.tcam_mask[2][440][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][441][0]=80'h0000000038f48a68b142;
sos_loop[0].somModel.tcam_mask[2][441][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][442][0]=80'h000000009759c188b4fd;
sos_loop[0].somModel.tcam_mask[2][442][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][443][0]=80'h00000000a08c0f3399b6;
sos_loop[0].somModel.tcam_mask[2][443][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][444][0]=80'h00000000820dea118ef9;
sos_loop[0].somModel.tcam_mask[2][444][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][445][0]=80'h00000000786f4fec3569;
sos_loop[0].somModel.tcam_mask[2][445][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][446][0]=80'h0000000035502a9bf339;
sos_loop[0].somModel.tcam_mask[2][446][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][447][0]=80'h00000000ede032f81911;
sos_loop[0].somModel.tcam_mask[2][447][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][448][0]=80'h00000000005d2da41d57;
sos_loop[0].somModel.tcam_mask[2][448][0]=80'hffffffffff8000000000;
sos_loop[0].somModel.tcam_data[2][449][0]=80'h000000001d551e45233a;
sos_loop[0].somModel.tcam_mask[2][449][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][450][0]=80'h000000001232e7e21619;
sos_loop[0].somModel.tcam_mask[2][450][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][451][0]=80'h000000009656bf8e0b9d;
sos_loop[0].somModel.tcam_mask[2][451][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][452][0]=80'h00000000282df63c9a42;
sos_loop[0].somModel.tcam_mask[2][452][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][453][0]=80'h00000000fb8cfa3efc1a;
sos_loop[0].somModel.tcam_mask[2][453][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][454][0]=80'h00000000e202a5e04142;
sos_loop[0].somModel.tcam_mask[2][454][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][455][0]=80'h00000000ce14bd93ed55;
sos_loop[0].somModel.tcam_mask[2][455][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][456][0]=80'h000000000b29b6b75332;
sos_loop[0].somModel.tcam_mask[2][456][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][457][0]=80'h00000000a560cfe7acfc;
sos_loop[0].somModel.tcam_mask[2][457][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][458][0]=80'h0000000099c7f0448e01;
sos_loop[0].somModel.tcam_mask[2][458][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][459][0]=80'h000000001dc007e9c85a;
sos_loop[0].somModel.tcam_mask[2][459][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][460][0]=80'h00000000d5bbfcebded1;
sos_loop[0].somModel.tcam_mask[2][460][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][461][0]=80'h000000007a59ce859cc7;
sos_loop[0].somModel.tcam_mask[2][461][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][462][0]=80'h000000004ea8c5b70bda;
sos_loop[0].somModel.tcam_mask[2][462][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][463][0]=80'h0000000052f1807fc08a;
sos_loop[0].somModel.tcam_mask[2][463][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][464][0]=80'h00000000206171d9529a;
sos_loop[0].somModel.tcam_mask[2][464][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][465][0]=80'h00000000498a7ea9d6a4;
sos_loop[0].somModel.tcam_mask[2][465][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][466][0]=80'h0000000068b1d8990008;
sos_loop[0].somModel.tcam_mask[2][466][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][467][0]=80'h00000000dfdd7f5c6649;
sos_loop[0].somModel.tcam_mask[2][467][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][468][0]=80'h00000000423c83f43d47;
sos_loop[0].somModel.tcam_mask[2][468][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][469][0]=80'h0000000071daa74440c3;
sos_loop[0].somModel.tcam_mask[2][469][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][470][0]=80'h000000006b7caeb2cb69;
sos_loop[0].somModel.tcam_mask[2][470][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][471][0]=80'h000000009301716b199f;
sos_loop[0].somModel.tcam_mask[2][471][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][472][0]=80'h00000000f30c2c261355;
sos_loop[0].somModel.tcam_mask[2][472][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][473][0]=80'h00000000e1037b5789b6;
sos_loop[0].somModel.tcam_mask[2][473][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][474][0]=80'h000000004ac85c163c30;
sos_loop[0].somModel.tcam_mask[2][474][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][475][0]=80'h00000000bd2e17a3bd71;
sos_loop[0].somModel.tcam_mask[2][475][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][476][0]=80'h000000008cfbaac12a25;
sos_loop[0].somModel.tcam_mask[2][476][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][477][0]=80'h00000000e07f86b355a4;
sos_loop[0].somModel.tcam_mask[2][477][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][478][0]=80'h00000000e24b3b5f435d;
sos_loop[0].somModel.tcam_mask[2][478][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][479][0]=80'h00000000c6100a3221e3;
sos_loop[0].somModel.tcam_mask[2][479][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][480][0]=80'h00000000d601e9e5d6ac;
sos_loop[0].somModel.tcam_mask[2][480][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][481][0]=80'h00000000a2ee82f9007b;
sos_loop[0].somModel.tcam_mask[2][481][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][482][0]=80'h00000000b4baf8944204;
sos_loop[0].somModel.tcam_mask[2][482][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][483][0]=80'h0000000078c5ee1f506d;
sos_loop[0].somModel.tcam_mask[2][483][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][484][0]=80'h0000000094176a64d950;
sos_loop[0].somModel.tcam_mask[2][484][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][485][0]=80'h00000000bdc7edf2bed3;
sos_loop[0].somModel.tcam_mask[2][485][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][486][0]=80'h00000000f6141087125a;
sos_loop[0].somModel.tcam_mask[2][486][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][487][0]=80'h000000004d8a6c4bb175;
sos_loop[0].somModel.tcam_mask[2][487][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][488][0]=80'h00000000d702b7ff755e;
sos_loop[0].somModel.tcam_mask[2][488][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][489][0]=80'h0000000017ad459c4491;
sos_loop[0].somModel.tcam_mask[2][489][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][490][0]=80'h00000000becd69de0af5;
sos_loop[0].somModel.tcam_mask[2][490][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][491][0]=80'h000000006db83a09cb40;
sos_loop[0].somModel.tcam_mask[2][491][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][492][0]=80'h00000000c15a3192c54e;
sos_loop[0].somModel.tcam_mask[2][492][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][493][0]=80'h00000000372729de79a7;
sos_loop[0].somModel.tcam_mask[2][493][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][494][0]=80'h00000000b7d5a573112e;
sos_loop[0].somModel.tcam_mask[2][494][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][495][0]=80'h00000000e7598a8d64ef;
sos_loop[0].somModel.tcam_mask[2][495][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][496][0]=80'h000000004d77a8f186e8;
sos_loop[0].somModel.tcam_mask[2][496][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][497][0]=80'h00000000b3a7e8c62438;
sos_loop[0].somModel.tcam_mask[2][497][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][498][0]=80'h000000005e628e40bad8;
sos_loop[0].somModel.tcam_mask[2][498][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][499][0]=80'h000000002c6ae9566a81;
sos_loop[0].somModel.tcam_mask[2][499][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][500][0]=80'h000000007c8088a4d780;
sos_loop[0].somModel.tcam_mask[2][500][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][501][0]=80'h00000000449da718991b;
sos_loop[0].somModel.tcam_mask[2][501][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][502][0]=80'h00000000eb14915c851e;
sos_loop[0].somModel.tcam_mask[2][502][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][503][0]=80'h000000003527b3d245b5;
sos_loop[0].somModel.tcam_mask[2][503][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][504][0]=80'h0000000085d7cc131a8a;
sos_loop[0].somModel.tcam_mask[2][504][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][505][0]=80'h00000000b448dcc734b3;
sos_loop[0].somModel.tcam_mask[2][505][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][506][0]=80'h000000000463282aaf56;
sos_loop[0].somModel.tcam_mask[2][506][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][507][0]=80'h00000000e6f6fe35b667;
sos_loop[0].somModel.tcam_mask[2][507][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][508][0]=80'h0000000080c258b15826;
sos_loop[0].somModel.tcam_mask[2][508][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][509][0]=80'h00000000faac4f7283f1;
sos_loop[0].somModel.tcam_mask[2][509][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][510][0]=80'h00000000a03cce697a88;
sos_loop[0].somModel.tcam_mask[2][510][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][511][0]=80'h00000000df03c7e186d0;
sos_loop[0].somModel.tcam_mask[2][511][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][512][0]=80'h00000000c301b2ddb491;
sos_loop[0].somModel.tcam_mask[2][512][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][513][0]=80'h0000000005a553a6d946;
sos_loop[0].somModel.tcam_mask[2][513][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][514][0]=80'h00000000ec81a0ecf565;
sos_loop[0].somModel.tcam_mask[2][514][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][515][0]=80'h0000000025b7ba6c7a22;
sos_loop[0].somModel.tcam_mask[2][515][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][516][0]=80'h00000000ff62f77af68e;
sos_loop[0].somModel.tcam_mask[2][516][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][517][0]=80'h0000000090696c0e7c49;
sos_loop[0].somModel.tcam_mask[2][517][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][518][0]=80'h00000000db542752b51b;
sos_loop[0].somModel.tcam_mask[2][518][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][519][0]=80'h000000005c669d7e5719;
sos_loop[0].somModel.tcam_mask[2][519][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][520][0]=80'h0000000007869b90d6d6;
sos_loop[0].somModel.tcam_mask[2][520][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][521][0]=80'h000000006ab3f4028bc4;
sos_loop[0].somModel.tcam_mask[2][521][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][522][0]=80'h00000000faf254c81784;
sos_loop[0].somModel.tcam_mask[2][522][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][523][0]=80'h00000000e91e80ddf2b6;
sos_loop[0].somModel.tcam_mask[2][523][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][524][0]=80'h0000000012ec8002dccf;
sos_loop[0].somModel.tcam_mask[2][524][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][525][0]=80'h000000001fb66119b301;
sos_loop[0].somModel.tcam_mask[2][525][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][526][0]=80'h0000000035cfa56dca6a;
sos_loop[0].somModel.tcam_mask[2][526][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][527][0]=80'h00000000257f17287640;
sos_loop[0].somModel.tcam_mask[2][527][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][528][0]=80'h00000000e24b719e5fd5;
sos_loop[0].somModel.tcam_mask[2][528][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][529][0]=80'h000000001b6de98d63bb;
sos_loop[0].somModel.tcam_mask[2][529][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][530][0]=80'h00000000c7396a1e1d0b;
sos_loop[0].somModel.tcam_mask[2][530][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][531][0]=80'h000000007fb43ae9cd4b;
sos_loop[0].somModel.tcam_mask[2][531][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][532][0]=80'h00000000a389a8825008;
sos_loop[0].somModel.tcam_mask[2][532][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][533][0]=80'h0000000062002cc089d3;
sos_loop[0].somModel.tcam_mask[2][533][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][534][0]=80'h00000000a2fc3e097fd8;
sos_loop[0].somModel.tcam_mask[2][534][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][535][0]=80'h0000000093938f2e7bb6;
sos_loop[0].somModel.tcam_mask[2][535][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][536][0]=80'h000000004c0878c8f3c9;
sos_loop[0].somModel.tcam_mask[2][536][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][537][0]=80'h000000006dad4681d74b;
sos_loop[0].somModel.tcam_mask[2][537][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][538][0]=80'h0000000090d849afd440;
sos_loop[0].somModel.tcam_mask[2][538][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][539][0]=80'h0000000099cea5c192b2;
sos_loop[0].somModel.tcam_mask[2][539][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][540][0]=80'h00000000439a63924ef9;
sos_loop[0].somModel.tcam_mask[2][540][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][541][0]=80'h0000000022efe4c3db4e;
sos_loop[0].somModel.tcam_mask[2][541][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][542][0]=80'h00000000935f8ae1eaca;
sos_loop[0].somModel.tcam_mask[2][542][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][543][0]=80'h00000000980ce89cb3ca;
sos_loop[0].somModel.tcam_mask[2][543][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][544][0]=80'h00000000b2b1d54e6143;
sos_loop[0].somModel.tcam_mask[2][544][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][545][0]=80'h00000000985262ca09c2;
sos_loop[0].somModel.tcam_mask[2][545][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][546][0]=80'h000000001b5370c23148;
sos_loop[0].somModel.tcam_mask[2][546][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][547][0]=80'h00000000fa6e44897737;
sos_loop[0].somModel.tcam_mask[2][547][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][548][0]=80'h00000000edc347b5f551;
sos_loop[0].somModel.tcam_mask[2][548][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][549][0]=80'h00000000bbafbcb86844;
sos_loop[0].somModel.tcam_mask[2][549][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][550][0]=80'h000000007fb9ba95cb59;
sos_loop[0].somModel.tcam_mask[2][550][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][551][0]=80'h00000000be931b35ee21;
sos_loop[0].somModel.tcam_mask[2][551][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][552][0]=80'h0000000039f56d709e34;
sos_loop[0].somModel.tcam_mask[2][552][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][553][0]=80'h000000004e9dfa08200a;
sos_loop[0].somModel.tcam_mask[2][553][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][554][0]=80'h00000000820c31b21a45;
sos_loop[0].somModel.tcam_mask[2][554][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][555][0]=80'h0000000005c7809f7005;
sos_loop[0].somModel.tcam_mask[2][555][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][556][0]=80'h000000003aca0c094cca;
sos_loop[0].somModel.tcam_mask[2][556][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][557][0]=80'h00000000745ae42f60b0;
sos_loop[0].somModel.tcam_mask[2][557][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][558][0]=80'h000000009ab1034e7c6e;
sos_loop[0].somModel.tcam_mask[2][558][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][559][0]=80'h000000008b03e00b02c2;
sos_loop[0].somModel.tcam_mask[2][559][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][560][0]=80'h00000000291393c268aa;
sos_loop[0].somModel.tcam_mask[2][560][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][561][0]=80'h000000004f5dda910b46;
sos_loop[0].somModel.tcam_mask[2][561][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][562][0]=80'h000000000d702572b740;
sos_loop[0].somModel.tcam_mask[2][562][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][563][0]=80'h0000000082eb751a50eb;
sos_loop[0].somModel.tcam_mask[2][563][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][564][0]=80'h0000000069f1bf212be5;
sos_loop[0].somModel.tcam_mask[2][564][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][565][0]=80'h00000000692f8eeae2e9;
sos_loop[0].somModel.tcam_mask[2][565][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][566][0]=80'h0000000019a683169415;
sos_loop[0].somModel.tcam_mask[2][566][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][567][0]=80'h0000000093bac3e6e685;
sos_loop[0].somModel.tcam_mask[2][567][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][568][0]=80'h000000004993bee769ac;
sos_loop[0].somModel.tcam_mask[2][568][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][569][0]=80'h00000000cd7fb4cb6753;
sos_loop[0].somModel.tcam_mask[2][569][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][570][0]=80'h000000000240e7a3c36d;
sos_loop[0].somModel.tcam_mask[2][570][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[2][571][0]=80'h00000000dee7cb29be85;
sos_loop[0].somModel.tcam_mask[2][571][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][572][0]=80'h00000000992597565e42;
sos_loop[0].somModel.tcam_mask[2][572][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][573][0]=80'h000000005cf48819c736;
sos_loop[0].somModel.tcam_mask[2][573][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][574][0]=80'h0000000047abe210da7f;
sos_loop[0].somModel.tcam_mask[2][574][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][575][0]=80'h00000000f93a1757baa0;
sos_loop[0].somModel.tcam_mask[2][575][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][576][0]=80'h000000007c1ceb4afc56;
sos_loop[0].somModel.tcam_mask[2][576][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][577][0]=80'h00000000af7d256d7cc4;
sos_loop[0].somModel.tcam_mask[2][577][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][578][0]=80'h0000000056f4eacb32c7;
sos_loop[0].somModel.tcam_mask[2][578][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][579][0]=80'h00000000b0d1add53e47;
sos_loop[0].somModel.tcam_mask[2][579][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][580][0]=80'h00000000d2755cc4bd17;
sos_loop[0].somModel.tcam_mask[2][580][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][581][0]=80'h00000000a6985589f9f2;
sos_loop[0].somModel.tcam_mask[2][581][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][582][0]=80'h00000000c617a79d7ece;
sos_loop[0].somModel.tcam_mask[2][582][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][583][0]=80'h00000000ce74602fffba;
sos_loop[0].somModel.tcam_mask[2][583][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][584][0]=80'h00000000f924b4b96d61;
sos_loop[0].somModel.tcam_mask[2][584][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][585][0]=80'h000000008c0b6b9901dc;
sos_loop[0].somModel.tcam_mask[2][585][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][586][0]=80'h00000000f68af87708bf;
sos_loop[0].somModel.tcam_mask[2][586][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][587][0]=80'h0000000074fa5f30fe3f;
sos_loop[0].somModel.tcam_mask[2][587][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][588][0]=80'h000000004db8a921b1d2;
sos_loop[0].somModel.tcam_mask[2][588][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][589][0]=80'h0000000018a72f979e24;
sos_loop[0].somModel.tcam_mask[2][589][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][590][0]=80'h00000000595e18260e26;
sos_loop[0].somModel.tcam_mask[2][590][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][591][0]=80'h00000000aad2d483e822;
sos_loop[0].somModel.tcam_mask[2][591][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][592][0]=80'h00000000343913fad305;
sos_loop[0].somModel.tcam_mask[2][592][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][593][0]=80'h00000000b3d2b6c10e97;
sos_loop[0].somModel.tcam_mask[2][593][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][594][0]=80'h000000005b359f4f70b0;
sos_loop[0].somModel.tcam_mask[2][594][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][595][0]=80'h00000000910fdf65238e;
sos_loop[0].somModel.tcam_mask[2][595][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][596][0]=80'h00000000858d2a03d342;
sos_loop[0].somModel.tcam_mask[2][596][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][597][0]=80'h0000000060c0b6079327;
sos_loop[0].somModel.tcam_mask[2][597][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][598][0]=80'h00000000ac7bf03559d7;
sos_loop[0].somModel.tcam_mask[2][598][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][599][0]=80'h000000009ad2390bbe32;
sos_loop[0].somModel.tcam_mask[2][599][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][600][0]=80'h00000000fa4f7ce06718;
sos_loop[0].somModel.tcam_mask[2][600][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][601][0]=80'h00000000d16fe65ec39f;
sos_loop[0].somModel.tcam_mask[2][601][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][602][0]=80'h000000002d99e55053a9;
sos_loop[0].somModel.tcam_mask[2][602][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][603][0]=80'h000000005159029f3697;
sos_loop[0].somModel.tcam_mask[2][603][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][604][0]=80'h00000000b4b0447b5549;
sos_loop[0].somModel.tcam_mask[2][604][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][605][0]=80'h00000000377b752a37b6;
sos_loop[0].somModel.tcam_mask[2][605][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][606][0]=80'h00000000220bb11437f4;
sos_loop[0].somModel.tcam_mask[2][606][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][607][0]=80'h00000000abd69fb1204e;
sos_loop[0].somModel.tcam_mask[2][607][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][608][0]=80'h00000000eb47988d0d8b;
sos_loop[0].somModel.tcam_mask[2][608][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][609][0]=80'h00000000ca9cc767edce;
sos_loop[0].somModel.tcam_mask[2][609][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][610][0]=80'h000000003b6f42cbe0a9;
sos_loop[0].somModel.tcam_mask[2][610][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][611][0]=80'h000000001dd3fa287076;
sos_loop[0].somModel.tcam_mask[2][611][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][612][0]=80'h000000009628912dbff2;
sos_loop[0].somModel.tcam_mask[2][612][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][613][0]=80'h0000000089a7951bea35;
sos_loop[0].somModel.tcam_mask[2][613][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][614][0]=80'h00000000c7b2ff90ab75;
sos_loop[0].somModel.tcam_mask[2][614][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][615][0]=80'h000000007ec37d3f35d1;
sos_loop[0].somModel.tcam_mask[2][615][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][616][0]=80'h00000000486d45350ba4;
sos_loop[0].somModel.tcam_mask[2][616][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][617][0]=80'h00000000f7c78a4aeffd;
sos_loop[0].somModel.tcam_mask[2][617][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][618][0]=80'h00000000ea7f3c4470a0;
sos_loop[0].somModel.tcam_mask[2][618][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][619][0]=80'h0000000095398bca46db;
sos_loop[0].somModel.tcam_mask[2][619][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][620][0]=80'h0000000002a21d269ef9;
sos_loop[0].somModel.tcam_mask[2][620][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[2][621][0]=80'h000000005ff142432afa;
sos_loop[0].somModel.tcam_mask[2][621][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][622][0]=80'h000000008d346fc65e2b;
sos_loop[0].somModel.tcam_mask[2][622][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][623][0]=80'h000000001a6584f50556;
sos_loop[0].somModel.tcam_mask[2][623][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][624][0]=80'h0000000008386da1029f;
sos_loop[0].somModel.tcam_mask[2][624][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][625][0]=80'h00000000db56c981ece6;
sos_loop[0].somModel.tcam_mask[2][625][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][626][0]=80'h00000000cfe8af38f522;
sos_loop[0].somModel.tcam_mask[2][626][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][627][0]=80'h000000008e919d8a745b;
sos_loop[0].somModel.tcam_mask[2][627][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][628][0]=80'h00000000543818958c78;
sos_loop[0].somModel.tcam_mask[2][628][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][629][0]=80'h00000000a8b931f97188;
sos_loop[0].somModel.tcam_mask[2][629][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][630][0]=80'h000000007dee0d849922;
sos_loop[0].somModel.tcam_mask[2][630][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][631][0]=80'h000000001017ca8a2953;
sos_loop[0].somModel.tcam_mask[2][631][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][632][0]=80'h000000007ed9cae24403;
sos_loop[0].somModel.tcam_mask[2][632][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][633][0]=80'h00000000ea187ed4d55a;
sos_loop[0].somModel.tcam_mask[2][633][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][634][0]=80'h000000002e76e28270f1;
sos_loop[0].somModel.tcam_mask[2][634][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][635][0]=80'h00000000f1980343333f;
sos_loop[0].somModel.tcam_mask[2][635][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][636][0]=80'h000000008de1c963c062;
sos_loop[0].somModel.tcam_mask[2][636][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][637][0]=80'h000000003fd86ea44501;
sos_loop[0].somModel.tcam_mask[2][637][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][638][0]=80'h00000000dc791a00bf2c;
sos_loop[0].somModel.tcam_mask[2][638][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][639][0]=80'h0000000076fd772b3105;
sos_loop[0].somModel.tcam_mask[2][639][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][640][0]=80'h000000009137a6d429b2;
sos_loop[0].somModel.tcam_mask[2][640][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][641][0]=80'h0000000049d4cbef7ccc;
sos_loop[0].somModel.tcam_mask[2][641][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][642][0]=80'h000000008051f12b529f;
sos_loop[0].somModel.tcam_mask[2][642][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][643][0]=80'h0000000008d6aa657a5e;
sos_loop[0].somModel.tcam_mask[2][643][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][644][0]=80'h0000000044bafb829ee6;
sos_loop[0].somModel.tcam_mask[2][644][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][645][0]=80'h00000000e55061ccc7b7;
sos_loop[0].somModel.tcam_mask[2][645][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][646][0]=80'h00000000d75970bd3bb0;
sos_loop[0].somModel.tcam_mask[2][646][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][647][0]=80'h000000004811729ba385;
sos_loop[0].somModel.tcam_mask[2][647][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][648][0]=80'h00000000c0501fd955df;
sos_loop[0].somModel.tcam_mask[2][648][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][649][0]=80'h00000000659c29b06d69;
sos_loop[0].somModel.tcam_mask[2][649][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][650][0]=80'h000000006aec373261a3;
sos_loop[0].somModel.tcam_mask[2][650][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][651][0]=80'h00000000c25cd90f5dab;
sos_loop[0].somModel.tcam_mask[2][651][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][652][0]=80'h00000000cee3230bfef6;
sos_loop[0].somModel.tcam_mask[2][652][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][653][0]=80'h000000007bde198a992f;
sos_loop[0].somModel.tcam_mask[2][653][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][654][0]=80'h000000007cd4d9587ccb;
sos_loop[0].somModel.tcam_mask[2][654][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][655][0]=80'h000000005cee7e94dd42;
sos_loop[0].somModel.tcam_mask[2][655][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][656][0]=80'h000000000c7f2c96b613;
sos_loop[0].somModel.tcam_mask[2][656][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][657][0]=80'h00000000f2de9d0bdde4;
sos_loop[0].somModel.tcam_mask[2][657][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][658][0]=80'h00000000b80342294761;
sos_loop[0].somModel.tcam_mask[2][658][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][659][0]=80'h00000000ef05f9051dde;
sos_loop[0].somModel.tcam_mask[2][659][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][660][0]=80'h00000000089d9864b0f7;
sos_loop[0].somModel.tcam_mask[2][660][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[2][661][0]=80'h00000000f84ebc6b5933;
sos_loop[0].somModel.tcam_mask[2][661][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][662][0]=80'h0000000099c7ebd6ef11;
sos_loop[0].somModel.tcam_mask[2][662][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][663][0]=80'h00000000a5cfc726453c;
sos_loop[0].somModel.tcam_mask[2][663][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][664][0]=80'h000000008e33ccc43905;
sos_loop[0].somModel.tcam_mask[2][664][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][665][0]=80'h0000000061dbc393f8b8;
sos_loop[0].somModel.tcam_mask[2][665][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][666][0]=80'h00000000b5776eb8e40c;
sos_loop[0].somModel.tcam_mask[2][666][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][667][0]=80'h00000000c56f02fbb8af;
sos_loop[0].somModel.tcam_mask[2][667][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][668][0]=80'h00000000f06ac89a6e2e;
sos_loop[0].somModel.tcam_mask[2][668][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][669][0]=80'h000000004d46ea5704c7;
sos_loop[0].somModel.tcam_mask[2][669][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][670][0]=80'h00000000018a0d2ab536;
sos_loop[0].somModel.tcam_mask[2][670][0]=80'hfffffffffe0000000000;
sos_loop[0].somModel.tcam_data[2][671][0]=80'h00000000de24ea9c8559;
sos_loop[0].somModel.tcam_mask[2][671][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][672][0]=80'h00000000117c2dcb8a3f;
sos_loop[0].somModel.tcam_mask[2][672][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][673][0]=80'h00000000042c5800a198;
sos_loop[0].somModel.tcam_mask[2][673][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][674][0]=80'h00000000c866641162c8;
sos_loop[0].somModel.tcam_mask[2][674][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][675][0]=80'h00000000c59ce2a178ef;
sos_loop[0].somModel.tcam_mask[2][675][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][676][0]=80'h0000000091b9a88b2186;
sos_loop[0].somModel.tcam_mask[2][676][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][677][0]=80'h00000000baaaa92f9330;
sos_loop[0].somModel.tcam_mask[2][677][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][678][0]=80'h00000000899bc4d45fed;
sos_loop[0].somModel.tcam_mask[2][678][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][679][0]=80'h0000000031aba86c07cd;
sos_loop[0].somModel.tcam_mask[2][679][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][680][0]=80'h00000000c4984e56b9a3;
sos_loop[0].somModel.tcam_mask[2][680][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][681][0]=80'h000000001b2cb5378bd2;
sos_loop[0].somModel.tcam_mask[2][681][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[2][682][0]=80'h00000000ff120ca68f9a;
sos_loop[0].somModel.tcam_mask[2][682][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][683][0]=80'h00000000a835dfd4a64e;
sos_loop[0].somModel.tcam_mask[2][683][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][684][0]=80'h00000000cc35683c57dc;
sos_loop[0].somModel.tcam_mask[2][684][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][685][0]=80'h00000000a5c1099a0ccc;
sos_loop[0].somModel.tcam_mask[2][685][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][686][0]=80'h00000000efd95c4e5fe9;
sos_loop[0].somModel.tcam_mask[2][686][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][687][0]=80'h000000007c76d25796aa;
sos_loop[0].somModel.tcam_mask[2][687][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][688][0]=80'h0000000007b60730923d;
sos_loop[0].somModel.tcam_mask[2][688][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][689][0]=80'h0000000007373b8b8f3c;
sos_loop[0].somModel.tcam_mask[2][689][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[2][690][0]=80'h0000000037e56c799b77;
sos_loop[0].somModel.tcam_mask[2][690][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[2][691][0]=80'h0000000064aeec7ab84c;
sos_loop[0].somModel.tcam_mask[2][691][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][692][0]=80'h00000000dc1814387312;
sos_loop[0].somModel.tcam_mask[2][692][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][693][0]=80'h00000000dd2835b8c4f9;
sos_loop[0].somModel.tcam_mask[2][693][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][694][0]=80'h000000005af2eb552cca;
sos_loop[0].somModel.tcam_mask[2][694][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][695][0]=80'h00000000446b9299fa74;
sos_loop[0].somModel.tcam_mask[2][695][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][696][0]=80'h0000000086928cf64fc6;
sos_loop[0].somModel.tcam_mask[2][696][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][697][0]=80'h00000000c4fdc019c61f;
sos_loop[0].somModel.tcam_mask[2][697][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][698][0]=80'h00000000882f97bb161f;
sos_loop[0].somModel.tcam_mask[2][698][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[2][699][0]=80'h000000004ed606f4518d;
sos_loop[0].somModel.tcam_mask[2][699][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[2][700][0]=80'h00000000bd46a3aa3c15;
sos_loop[0].somModel.tcam_mask[2][700][0]=80'hffffffff000000000000;
sos_loop[0].somModel.sram_dat[2][0][0]=96'hdeadbf;
sos_loop[0].somModel.sram_ptr[2][0]=939;
sos_loop[0].somModel.sram_dat[2][1][0]=96'h7f1ea9;
sos_loop[0].somModel.sram_ptr[2][1]=2;
sos_loop[0].somModel.sram_dat[2][2][0]=96'h18d7d4;
sos_loop[0].somModel.sram_ptr[2][2]=2;
sos_loop[0].somModel.sram_dat[2][3][0]=96'h879503;
sos_loop[0].somModel.sram_ptr[2][3]=2;
sos_loop[0].somModel.sram_dat[2][4][0]=96'h795e9d;
sos_loop[0].somModel.sram_ptr[2][4]=2;
sos_loop[0].somModel.sram_dat[2][5][0]=96'hd8811f;
sos_loop[0].somModel.sram_ptr[2][5]=2;
sos_loop[0].somModel.sram_dat[2][6][0]=96'hf72c4f;
sos_loop[0].somModel.sram_ptr[2][6]=2;
sos_loop[0].somModel.sram_dat[2][7][0]=96'h45bc37;
sos_loop[0].somModel.sram_ptr[2][7]=2;
sos_loop[0].somModel.sram_dat[2][8][0]=96'ha9ca1e;
sos_loop[0].somModel.sram_ptr[2][8]=2;
sos_loop[0].somModel.sram_dat[2][9][0]=96'h95fadc;
sos_loop[0].somModel.sram_ptr[2][9]=2;
sos_loop[0].somModel.sram_dat[2][10][0]=96'hfd7856;
sos_loop[0].somModel.sram_ptr[2][10]=2;
sos_loop[0].somModel.sram_dat[2][11][0]=96'h3ac1d0;
sos_loop[0].somModel.sram_ptr[2][11]=2;
sos_loop[0].somModel.sram_dat[2][12][0]=96'hc47e0;
sos_loop[0].somModel.sram_ptr[2][12]=2;
sos_loop[0].somModel.sram_dat[2][13][0]=96'hfb27f9;
sos_loop[0].somModel.sram_ptr[2][13]=2;
sos_loop[0].somModel.sram_dat[2][14][0]=96'h18fca4;
sos_loop[0].somModel.sram_ptr[2][14]=2;
sos_loop[0].somModel.sram_dat[2][15][0]=96'h2e4356;
sos_loop[0].somModel.sram_ptr[2][15]=2;
sos_loop[0].somModel.sram_dat[2][16][0]=96'h56a40c;
sos_loop[0].somModel.sram_ptr[2][16]=2;
sos_loop[0].somModel.sram_dat[2][17][0]=96'h18540e;
sos_loop[0].somModel.sram_ptr[2][17]=2;
sos_loop[0].somModel.sram_dat[2][18][0]=96'hea2b44;
sos_loop[0].somModel.sram_ptr[2][18]=2;
sos_loop[0].somModel.sram_dat[2][19][0]=96'h84c769;
sos_loop[0].somModel.sram_ptr[2][19]=2;
sos_loop[0].somModel.sram_dat[2][20][0]=96'h9ae0b9;
sos_loop[0].somModel.sram_ptr[2][20]=2;
sos_loop[0].somModel.sram_dat[2][21][0]=96'ha15356;
sos_loop[0].somModel.sram_ptr[2][21]=2;
sos_loop[0].somModel.sram_dat[2][22][0]=96'h5a0605;
sos_loop[0].somModel.sram_ptr[2][22]=2;
sos_loop[0].somModel.sram_dat[2][23][0]=96'h6fe0cb;
sos_loop[0].somModel.sram_ptr[2][23]=2;
sos_loop[0].somModel.sram_dat[2][24][0]=96'he646d6;
sos_loop[0].somModel.sram_ptr[2][24]=2;
sos_loop[0].somModel.sram_dat[2][25][0]=96'ha2d6b;
sos_loop[0].somModel.sram_ptr[2][25]=2;
sos_loop[0].somModel.sram_dat[2][26][0]=96'hf04d5b;
sos_loop[0].somModel.sram_ptr[2][26]=2;
sos_loop[0].somModel.sram_dat[2][27][0]=96'h4c578c;
sos_loop[0].somModel.sram_ptr[2][27]=2;
sos_loop[0].somModel.sram_dat[2][28][0]=96'h888d1f;
sos_loop[0].somModel.sram_ptr[2][28]=2;
sos_loop[0].somModel.sram_dat[2][29][0]=96'h2ca3fe;
sos_loop[0].somModel.sram_ptr[2][29]=2;
sos_loop[0].somModel.sram_dat[2][30][0]=96'h63455b;
sos_loop[0].somModel.sram_ptr[2][30]=2;
sos_loop[0].somModel.sram_dat[2][31][0]=96'h2768c3;
sos_loop[0].somModel.sram_ptr[2][31]=2;
sos_loop[0].somModel.sram_dat[2][32][0]=96'h7cb8cb;
sos_loop[0].somModel.sram_ptr[2][32]=2;
sos_loop[0].somModel.sram_dat[2][33][0]=96'h62f735;
sos_loop[0].somModel.sram_ptr[2][33]=2;
sos_loop[0].somModel.sram_dat[2][34][0]=96'h2fa2ac;
sos_loop[0].somModel.sram_ptr[2][34]=2;
sos_loop[0].somModel.sram_dat[2][35][0]=96'h6b0b30;
sos_loop[0].somModel.sram_ptr[2][35]=2;
sos_loop[0].somModel.sram_dat[2][36][0]=96'hdc4120;
sos_loop[0].somModel.sram_ptr[2][36]=2;
sos_loop[0].somModel.sram_dat[2][37][0]=96'hd471aa;
sos_loop[0].somModel.sram_ptr[2][37]=2;
sos_loop[0].somModel.sram_dat[2][38][0]=96'h40a7fc;
sos_loop[0].somModel.sram_ptr[2][38]=2;
sos_loop[0].somModel.sram_dat[2][39][0]=96'hac33c6;
sos_loop[0].somModel.sram_ptr[2][39]=2;
sos_loop[0].somModel.sram_dat[2][40][0]=96'h109775;
sos_loop[0].somModel.sram_ptr[2][40]=2;
sos_loop[0].somModel.sram_dat[2][41][0]=96'hc3ff40;
sos_loop[0].somModel.sram_ptr[2][41]=2;
sos_loop[0].somModel.sram_dat[2][42][0]=96'h283e24;
sos_loop[0].somModel.sram_ptr[2][42]=2;
sos_loop[0].somModel.sram_dat[2][43][0]=96'hd2bca2;
sos_loop[0].somModel.sram_ptr[2][43]=2;
sos_loop[0].somModel.sram_dat[2][44][0]=96'h5178a5;
sos_loop[0].somModel.sram_ptr[2][44]=2;
sos_loop[0].somModel.sram_dat[2][45][0]=96'h9ab1a5;
sos_loop[0].somModel.sram_ptr[2][45]=2;
sos_loop[0].somModel.sram_dat[2][46][0]=96'hdd0418;
sos_loop[0].somModel.sram_ptr[2][46]=2;
sos_loop[0].somModel.sram_dat[2][47][0]=96'h4341e8;
sos_loop[0].somModel.sram_ptr[2][47]=2;
sos_loop[0].somModel.sram_dat[2][48][0]=96'hbeafd2;
sos_loop[0].somModel.sram_ptr[2][48]=2;
sos_loop[0].somModel.sram_dat[2][49][0]=96'h653c68;
sos_loop[0].somModel.sram_ptr[2][49]=2;
sos_loop[0].somModel.sram_dat[2][50][0]=96'hc2f7fb;
sos_loop[0].somModel.sram_ptr[2][50]=2;
sos_loop[0].somModel.sram_dat[2][51][0]=96'h2ec425;
sos_loop[0].somModel.sram_ptr[2][51]=2;
sos_loop[0].somModel.sram_dat[2][52][0]=96'h39f1b8;
sos_loop[0].somModel.sram_ptr[2][52]=2;
sos_loop[0].somModel.sram_dat[2][53][0]=96'h65b81f;
sos_loop[0].somModel.sram_ptr[2][53]=2;
sos_loop[0].somModel.sram_dat[2][54][0]=96'he84bff;
sos_loop[0].somModel.sram_ptr[2][54]=2;
sos_loop[0].somModel.sram_dat[2][55][0]=96'h6f12c1;
sos_loop[0].somModel.sram_ptr[2][55]=2;
sos_loop[0].somModel.sram_dat[2][56][0]=96'h638539;
sos_loop[0].somModel.sram_ptr[2][56]=2;
sos_loop[0].somModel.sram_dat[2][57][0]=96'h74386b;
sos_loop[0].somModel.sram_ptr[2][57]=2;
sos_loop[0].somModel.sram_dat[2][58][0]=96'h6ec296;
sos_loop[0].somModel.sram_ptr[2][58]=2;
sos_loop[0].somModel.sram_dat[2][59][0]=96'h9dc45a;
sos_loop[0].somModel.sram_ptr[2][59]=2;
sos_loop[0].somModel.sram_dat[2][60][0]=96'h7bdeb2;
sos_loop[0].somModel.sram_ptr[2][60]=2;
sos_loop[0].somModel.sram_dat[2][61][0]=96'h109400;
sos_loop[0].somModel.sram_ptr[2][61]=2;
sos_loop[0].somModel.sram_dat[2][62][0]=96'h3ed34b;
sos_loop[0].somModel.sram_ptr[2][62]=2;
sos_loop[0].somModel.sram_dat[2][63][0]=96'h83a39a;
sos_loop[0].somModel.sram_ptr[2][63]=2;
sos_loop[0].somModel.sram_dat[2][64][0]=96'hb39350;
sos_loop[0].somModel.sram_ptr[2][64]=2;
sos_loop[0].somModel.sram_dat[2][65][0]=96'h3fd68e;
sos_loop[0].somModel.sram_ptr[2][65]=2;
sos_loop[0].somModel.sram_dat[2][66][0]=96'h168dc8;
sos_loop[0].somModel.sram_ptr[2][66]=2;
sos_loop[0].somModel.sram_dat[2][67][0]=96'hc7d864;
sos_loop[0].somModel.sram_ptr[2][67]=2;
sos_loop[0].somModel.sram_dat[2][68][0]=96'h6ac4b8;
sos_loop[0].somModel.sram_ptr[2][68]=2;
sos_loop[0].somModel.sram_dat[2][69][0]=96'h29c5fa;
sos_loop[0].somModel.sram_ptr[2][69]=2;
sos_loop[0].somModel.sram_dat[2][70][0]=96'h7775e4;
sos_loop[0].somModel.sram_ptr[2][70]=2;
sos_loop[0].somModel.sram_dat[2][71][0]=96'h354a38;
sos_loop[0].somModel.sram_ptr[2][71]=2;
sos_loop[0].somModel.sram_dat[2][72][0]=96'h482f82;
sos_loop[0].somModel.sram_ptr[2][72]=2;
sos_loop[0].somModel.sram_dat[2][73][0]=96'h8f4dc7;
sos_loop[0].somModel.sram_ptr[2][73]=2;
sos_loop[0].somModel.sram_dat[2][74][0]=96'h2f794e;
sos_loop[0].somModel.sram_ptr[2][74]=2;
sos_loop[0].somModel.sram_dat[2][75][0]=96'hc688bd;
sos_loop[0].somModel.sram_ptr[2][75]=2;
sos_loop[0].somModel.sram_dat[2][76][0]=96'h8c6bf8;
sos_loop[0].somModel.sram_ptr[2][76]=2;
sos_loop[0].somModel.sram_dat[2][77][0]=96'h4a580d;
sos_loop[0].somModel.sram_ptr[2][77]=2;
sos_loop[0].somModel.sram_dat[2][78][0]=96'he51d07;
sos_loop[0].somModel.sram_ptr[2][78]=2;
sos_loop[0].somModel.sram_dat[2][79][0]=96'h6576cb;
sos_loop[0].somModel.sram_ptr[2][79]=2;
sos_loop[0].somModel.sram_dat[2][80][0]=96'h672b33;
sos_loop[0].somModel.sram_ptr[2][80]=2;
sos_loop[0].somModel.sram_dat[2][81][0]=96'h765369;
sos_loop[0].somModel.sram_ptr[2][81]=2;
sos_loop[0].somModel.sram_dat[2][82][0]=96'h65548;
sos_loop[0].somModel.sram_ptr[2][82]=2;
sos_loop[0].somModel.sram_dat[2][83][0]=96'hfa8b7f;
sos_loop[0].somModel.sram_ptr[2][83]=2;
sos_loop[0].somModel.sram_dat[2][84][0]=96'h9e0149;
sos_loop[0].somModel.sram_ptr[2][84]=2;
sos_loop[0].somModel.sram_dat[2][85][0]=96'h3700bc;
sos_loop[0].somModel.sram_ptr[2][85]=2;
sos_loop[0].somModel.sram_dat[2][86][0]=96'ha26d54;
sos_loop[0].somModel.sram_ptr[2][86]=2;
sos_loop[0].somModel.sram_dat[2][87][0]=96'h485e50;
sos_loop[0].somModel.sram_ptr[2][87]=2;
sos_loop[0].somModel.sram_dat[2][88][0]=96'h4e377c;
sos_loop[0].somModel.sram_ptr[2][88]=2;
sos_loop[0].somModel.sram_dat[2][89][0]=96'h290bd8;
sos_loop[0].somModel.sram_ptr[2][89]=2;
sos_loop[0].somModel.sram_dat[2][90][0]=96'h79eac3;
sos_loop[0].somModel.sram_ptr[2][90]=2;
sos_loop[0].somModel.sram_dat[2][91][0]=96'haeb963;
sos_loop[0].somModel.sram_ptr[2][91]=2;
sos_loop[0].somModel.sram_dat[2][92][0]=96'he60f6;
sos_loop[0].somModel.sram_ptr[2][92]=2;
sos_loop[0].somModel.sram_dat[2][93][0]=96'hebc64c;
sos_loop[0].somModel.sram_ptr[2][93]=2;
sos_loop[0].somModel.sram_dat[2][94][0]=96'hfd79da;
sos_loop[0].somModel.sram_ptr[2][94]=2;
sos_loop[0].somModel.sram_dat[2][95][0]=96'h5f903f;
sos_loop[0].somModel.sram_ptr[2][95]=2;
sos_loop[0].somModel.sram_dat[2][96][0]=96'h8c6098;
sos_loop[0].somModel.sram_ptr[2][96]=2;
sos_loop[0].somModel.sram_dat[2][97][0]=96'h52bbf8;
sos_loop[0].somModel.sram_ptr[2][97]=2;
sos_loop[0].somModel.sram_dat[2][98][0]=96'h67064a;
sos_loop[0].somModel.sram_ptr[2][98]=2;
sos_loop[0].somModel.sram_dat[2][99][0]=96'heda0ac;
sos_loop[0].somModel.sram_ptr[2][99]=2;
sos_loop[0].somModel.sram_dat[2][100][0]=96'h9fe0b2;
sos_loop[0].somModel.sram_ptr[2][100]=2;
sos_loop[0].somModel.sram_dat[2][101][0]=96'h2b0b9e;
sos_loop[0].somModel.sram_ptr[2][101]=2;
sos_loop[0].somModel.sram_dat[2][102][0]=96'h8ed315;
sos_loop[0].somModel.sram_ptr[2][102]=2;
sos_loop[0].somModel.sram_dat[2][103][0]=96'h3fa5eb;
sos_loop[0].somModel.sram_ptr[2][103]=2;
sos_loop[0].somModel.sram_dat[2][104][0]=96'hd5a9ea;
sos_loop[0].somModel.sram_ptr[2][104]=2;
sos_loop[0].somModel.sram_dat[2][105][0]=96'h3b5063;
sos_loop[0].somModel.sram_ptr[2][105]=2;
sos_loop[0].somModel.sram_dat[2][106][0]=96'h3de498;
sos_loop[0].somModel.sram_ptr[2][106]=2;
sos_loop[0].somModel.sram_dat[2][107][0]=96'h34d05b;
sos_loop[0].somModel.sram_ptr[2][107]=2;
sos_loop[0].somModel.sram_dat[2][108][0]=96'h9906b4;
sos_loop[0].somModel.sram_ptr[2][108]=2;
sos_loop[0].somModel.sram_dat[2][109][0]=96'h8e8559;
sos_loop[0].somModel.sram_ptr[2][109]=2;
sos_loop[0].somModel.sram_dat[2][110][0]=96'he3f52;
sos_loop[0].somModel.sram_ptr[2][110]=2;
sos_loop[0].somModel.sram_dat[2][111][0]=96'h4b4571;
sos_loop[0].somModel.sram_ptr[2][111]=2;
sos_loop[0].somModel.sram_dat[2][112][0]=96'h1da95e;
sos_loop[0].somModel.sram_ptr[2][112]=2;
sos_loop[0].somModel.sram_dat[2][113][0]=96'hf8a77d;
sos_loop[0].somModel.sram_ptr[2][113]=2;
sos_loop[0].somModel.sram_dat[2][114][0]=96'h773e7;
sos_loop[0].somModel.sram_ptr[2][114]=2;
sos_loop[0].somModel.sram_dat[2][115][0]=96'hcc18d8;
sos_loop[0].somModel.sram_ptr[2][115]=2;
sos_loop[0].somModel.sram_dat[2][116][0]=96'h523f2c;
sos_loop[0].somModel.sram_ptr[2][116]=2;
sos_loop[0].somModel.sram_dat[2][117][0]=96'hd32eb1;
sos_loop[0].somModel.sram_ptr[2][117]=2;
sos_loop[0].somModel.sram_dat[2][118][0]=96'hb10a04;
sos_loop[0].somModel.sram_ptr[2][118]=2;
sos_loop[0].somModel.sram_dat[2][119][0]=96'h9e289a;
sos_loop[0].somModel.sram_ptr[2][119]=2;
sos_loop[0].somModel.sram_dat[2][120][0]=96'h3f745c;
sos_loop[0].somModel.sram_ptr[2][120]=2;
sos_loop[0].somModel.sram_dat[2][121][0]=96'hb4d716;
sos_loop[0].somModel.sram_ptr[2][121]=2;
sos_loop[0].somModel.sram_dat[2][122][0]=96'h353aba;
sos_loop[0].somModel.sram_ptr[2][122]=2;
sos_loop[0].somModel.sram_dat[2][123][0]=96'h138266;
sos_loop[0].somModel.sram_ptr[2][123]=2;
sos_loop[0].somModel.sram_dat[2][124][0]=96'h98c3a8;
sos_loop[0].somModel.sram_ptr[2][124]=2;
sos_loop[0].somModel.sram_dat[2][125][0]=96'ha72bb0;
sos_loop[0].somModel.sram_ptr[2][125]=2;
sos_loop[0].somModel.sram_dat[2][126][0]=96'hf0a808;
sos_loop[0].somModel.sram_ptr[2][126]=2;
sos_loop[0].somModel.sram_dat[2][127][0]=96'h2ecc7c;
sos_loop[0].somModel.sram_ptr[2][127]=2;
sos_loop[0].somModel.sram_dat[2][128][0]=96'h70432e;
sos_loop[0].somModel.sram_ptr[2][128]=2;
sos_loop[0].somModel.sram_dat[2][129][0]=96'h9e5629;
sos_loop[0].somModel.sram_ptr[2][129]=2;
sos_loop[0].somModel.sram_dat[2][130][0]=96'hb9028f;
sos_loop[0].somModel.sram_ptr[2][130]=2;
sos_loop[0].somModel.sram_dat[2][131][0]=96'h7d192f;
sos_loop[0].somModel.sram_ptr[2][131]=2;
sos_loop[0].somModel.sram_dat[2][132][0]=96'h9f9291;
sos_loop[0].somModel.sram_ptr[2][132]=2;
sos_loop[0].somModel.sram_dat[2][133][0]=96'hee6a20;
sos_loop[0].somModel.sram_ptr[2][133]=2;
sos_loop[0].somModel.sram_dat[2][134][0]=96'h53672d;
sos_loop[0].somModel.sram_ptr[2][134]=2;
sos_loop[0].somModel.sram_dat[2][135][0]=96'hdd027c;
sos_loop[0].somModel.sram_ptr[2][135]=2;
sos_loop[0].somModel.sram_dat[2][136][0]=96'hdc08c;
sos_loop[0].somModel.sram_ptr[2][136]=2;
sos_loop[0].somModel.sram_dat[2][137][0]=96'h58402c;
sos_loop[0].somModel.sram_ptr[2][137]=2;
sos_loop[0].somModel.sram_dat[2][138][0]=96'hc81a4a;
sos_loop[0].somModel.sram_ptr[2][138]=2;
sos_loop[0].somModel.sram_dat[2][139][0]=96'hedd5d3;
sos_loop[0].somModel.sram_ptr[2][139]=2;
sos_loop[0].somModel.sram_dat[2][140][0]=96'h4b52;
sos_loop[0].somModel.sram_ptr[2][140]=2;
sos_loop[0].somModel.sram_dat[2][141][0]=96'he03ed4;
sos_loop[0].somModel.sram_ptr[2][141]=2;
sos_loop[0].somModel.sram_dat[2][142][0]=96'h7e9436;
sos_loop[0].somModel.sram_ptr[2][142]=2;
sos_loop[0].somModel.sram_dat[2][143][0]=96'h784bef;
sos_loop[0].somModel.sram_ptr[2][143]=2;
sos_loop[0].somModel.sram_dat[2][144][0]=96'h42f39d;
sos_loop[0].somModel.sram_ptr[2][144]=2;
sos_loop[0].somModel.sram_dat[2][145][0]=96'hbe6a7e;
sos_loop[0].somModel.sram_ptr[2][145]=2;
sos_loop[0].somModel.sram_dat[2][146][0]=96'h826f57;
sos_loop[0].somModel.sram_ptr[2][146]=2;
sos_loop[0].somModel.sram_dat[2][147][0]=96'h29e2c;
sos_loop[0].somModel.sram_ptr[2][147]=2;
sos_loop[0].somModel.sram_dat[2][148][0]=96'h29c960;
sos_loop[0].somModel.sram_ptr[2][148]=2;
sos_loop[0].somModel.sram_dat[2][149][0]=96'h19c756;
sos_loop[0].somModel.sram_ptr[2][149]=2;
sos_loop[0].somModel.sram_dat[2][150][0]=96'h1fbdf;
sos_loop[0].somModel.sram_ptr[2][150]=2;
sos_loop[0].somModel.sram_dat[2][151][0]=96'h798a3;
sos_loop[0].somModel.sram_ptr[2][151]=2;
sos_loop[0].somModel.sram_dat[2][152][0]=96'h376c99;
sos_loop[0].somModel.sram_ptr[2][152]=2;
sos_loop[0].somModel.sram_dat[2][153][0]=96'h2e7c93;
sos_loop[0].somModel.sram_ptr[2][153]=2;
sos_loop[0].somModel.sram_dat[2][154][0]=96'h6e0c48;
sos_loop[0].somModel.sram_ptr[2][154]=2;
sos_loop[0].somModel.sram_dat[2][155][0]=96'h7848e4;
sos_loop[0].somModel.sram_ptr[2][155]=2;
sos_loop[0].somModel.sram_dat[2][156][0]=96'heab49b;
sos_loop[0].somModel.sram_ptr[2][156]=2;
sos_loop[0].somModel.sram_dat[2][157][0]=96'h3c4183;
sos_loop[0].somModel.sram_ptr[2][157]=2;
sos_loop[0].somModel.sram_dat[2][158][0]=96'h206e77;
sos_loop[0].somModel.sram_ptr[2][158]=2;
sos_loop[0].somModel.sram_dat[2][159][0]=96'h60af7b;
sos_loop[0].somModel.sram_ptr[2][159]=2;
sos_loop[0].somModel.sram_dat[2][160][0]=96'h532847;
sos_loop[0].somModel.sram_ptr[2][160]=2;
sos_loop[0].somModel.sram_dat[2][161][0]=96'hbad608;
sos_loop[0].somModel.sram_ptr[2][161]=2;
sos_loop[0].somModel.sram_dat[2][162][0]=96'h47a19a;
sos_loop[0].somModel.sram_ptr[2][162]=2;
sos_loop[0].somModel.sram_dat[2][163][0]=96'hf8c422;
sos_loop[0].somModel.sram_ptr[2][163]=2;
sos_loop[0].somModel.sram_dat[2][164][0]=96'h9c50ab;
sos_loop[0].somModel.sram_ptr[2][164]=2;
sos_loop[0].somModel.sram_dat[2][165][0]=96'h2c4a16;
sos_loop[0].somModel.sram_ptr[2][165]=2;
sos_loop[0].somModel.sram_dat[2][166][0]=96'he2f212;
sos_loop[0].somModel.sram_ptr[2][166]=2;
sos_loop[0].somModel.sram_dat[2][167][0]=96'h32b6e2;
sos_loop[0].somModel.sram_ptr[2][167]=2;
sos_loop[0].somModel.sram_dat[2][168][0]=96'h501cd9;
sos_loop[0].somModel.sram_ptr[2][168]=2;
sos_loop[0].somModel.sram_dat[2][169][0]=96'h59d817;
sos_loop[0].somModel.sram_ptr[2][169]=2;
sos_loop[0].somModel.sram_dat[2][170][0]=96'h79c4b3;
sos_loop[0].somModel.sram_ptr[2][170]=2;
sos_loop[0].somModel.sram_dat[2][171][0]=96'hdbfb38;
sos_loop[0].somModel.sram_ptr[2][171]=2;
sos_loop[0].somModel.sram_dat[2][172][0]=96'h3c8d91;
sos_loop[0].somModel.sram_ptr[2][172]=2;
sos_loop[0].somModel.sram_dat[2][173][0]=96'h700b97;
sos_loop[0].somModel.sram_ptr[2][173]=2;
sos_loop[0].somModel.sram_dat[2][174][0]=96'h6a6798;
sos_loop[0].somModel.sram_ptr[2][174]=2;
sos_loop[0].somModel.sram_dat[2][175][0]=96'hb16541;
sos_loop[0].somModel.sram_ptr[2][175]=2;
sos_loop[0].somModel.sram_dat[2][176][0]=96'h148fdc;
sos_loop[0].somModel.sram_ptr[2][176]=2;
sos_loop[0].somModel.sram_dat[2][177][0]=96'hc77ae0;
sos_loop[0].somModel.sram_ptr[2][177]=2;
sos_loop[0].somModel.sram_dat[2][178][0]=96'h289a41;
sos_loop[0].somModel.sram_ptr[2][178]=2;
sos_loop[0].somModel.sram_dat[2][179][0]=96'hcce9c6;
sos_loop[0].somModel.sram_ptr[2][179]=2;
sos_loop[0].somModel.sram_dat[2][180][0]=96'h3293d0;
sos_loop[0].somModel.sram_ptr[2][180]=2;
sos_loop[0].somModel.sram_dat[2][181][0]=96'h85fe27;
sos_loop[0].somModel.sram_ptr[2][181]=2;
sos_loop[0].somModel.sram_dat[2][182][0]=96'h7de321;
sos_loop[0].somModel.sram_ptr[2][182]=2;
sos_loop[0].somModel.sram_dat[2][183][0]=96'h556878;
sos_loop[0].somModel.sram_ptr[2][183]=2;
sos_loop[0].somModel.sram_dat[2][184][0]=96'ha2e200;
sos_loop[0].somModel.sram_ptr[2][184]=2;
sos_loop[0].somModel.sram_dat[2][185][0]=96'hf7b199;
sos_loop[0].somModel.sram_ptr[2][185]=2;
sos_loop[0].somModel.sram_dat[2][186][0]=96'h4e7d0f;
sos_loop[0].somModel.sram_ptr[2][186]=2;
sos_loop[0].somModel.sram_dat[2][187][0]=96'h2932d5;
sos_loop[0].somModel.sram_ptr[2][187]=2;
sos_loop[0].somModel.sram_dat[2][188][0]=96'hf10ee2;
sos_loop[0].somModel.sram_ptr[2][188]=2;
sos_loop[0].somModel.sram_dat[2][189][0]=96'hd3cb30;
sos_loop[0].somModel.sram_ptr[2][189]=2;
sos_loop[0].somModel.sram_dat[2][190][0]=96'hdc4082;
sos_loop[0].somModel.sram_ptr[2][190]=2;
sos_loop[0].somModel.sram_dat[2][191][0]=96'h4680df;
sos_loop[0].somModel.sram_ptr[2][191]=2;
sos_loop[0].somModel.sram_dat[2][192][0]=96'h3e3ace;
sos_loop[0].somModel.sram_ptr[2][192]=2;
sos_loop[0].somModel.sram_dat[2][193][0]=96'h278237;
sos_loop[0].somModel.sram_ptr[2][193]=2;
sos_loop[0].somModel.sram_dat[2][194][0]=96'hf58b4b;
sos_loop[0].somModel.sram_ptr[2][194]=2;
sos_loop[0].somModel.sram_dat[2][195][0]=96'h53a60b;
sos_loop[0].somModel.sram_ptr[2][195]=2;
sos_loop[0].somModel.sram_dat[2][196][0]=96'h29bce4;
sos_loop[0].somModel.sram_ptr[2][196]=2;
sos_loop[0].somModel.sram_dat[2][197][0]=96'hbf1a0a;
sos_loop[0].somModel.sram_ptr[2][197]=2;
sos_loop[0].somModel.sram_dat[2][198][0]=96'he19318;
sos_loop[0].somModel.sram_ptr[2][198]=2;
sos_loop[0].somModel.sram_dat[2][199][0]=96'h44d266;
sos_loop[0].somModel.sram_ptr[2][199]=2;
sos_loop[0].somModel.sram_dat[2][200][0]=96'ha6b455;
sos_loop[0].somModel.sram_ptr[2][200]=2;
sos_loop[0].somModel.sram_dat[2][201][0]=96'ha1ed9d;
sos_loop[0].somModel.sram_ptr[2][201]=2;
sos_loop[0].somModel.sram_dat[2][202][0]=96'h4fc0f7;
sos_loop[0].somModel.sram_ptr[2][202]=2;
sos_loop[0].somModel.sram_dat[2][203][0]=96'h83eaaf;
sos_loop[0].somModel.sram_ptr[2][203]=2;
sos_loop[0].somModel.sram_dat[2][204][0]=96'h1d8f2;
sos_loop[0].somModel.sram_ptr[2][204]=2;
sos_loop[0].somModel.sram_dat[2][205][0]=96'hc8461;
sos_loop[0].somModel.sram_ptr[2][205]=2;
sos_loop[0].somModel.sram_dat[2][206][0]=96'h5a9ad8;
sos_loop[0].somModel.sram_ptr[2][206]=2;
sos_loop[0].somModel.sram_dat[2][207][0]=96'h45adc4;
sos_loop[0].somModel.sram_ptr[2][207]=2;
sos_loop[0].somModel.sram_dat[2][208][0]=96'h44e7f5;
sos_loop[0].somModel.sram_ptr[2][208]=2;
sos_loop[0].somModel.sram_dat[2][209][0]=96'h4a5dba;
sos_loop[0].somModel.sram_ptr[2][209]=2;
sos_loop[0].somModel.sram_dat[2][210][0]=96'h82d37a;
sos_loop[0].somModel.sram_ptr[2][210]=2;
sos_loop[0].somModel.sram_dat[2][211][0]=96'ha5936e;
sos_loop[0].somModel.sram_ptr[2][211]=2;
sos_loop[0].somModel.sram_dat[2][212][0]=96'h7b239;
sos_loop[0].somModel.sram_ptr[2][212]=2;
sos_loop[0].somModel.sram_dat[2][213][0]=96'h12fd45;
sos_loop[0].somModel.sram_ptr[2][213]=2;
sos_loop[0].somModel.sram_dat[2][214][0]=96'h842ec1;
sos_loop[0].somModel.sram_ptr[2][214]=2;
sos_loop[0].somModel.sram_dat[2][215][0]=96'h5fee07;
sos_loop[0].somModel.sram_ptr[2][215]=2;
sos_loop[0].somModel.sram_dat[2][216][0]=96'h386dc0;
sos_loop[0].somModel.sram_ptr[2][216]=2;
sos_loop[0].somModel.sram_dat[2][217][0]=96'h30a003;
sos_loop[0].somModel.sram_ptr[2][217]=2;
sos_loop[0].somModel.sram_dat[2][218][0]=96'h69dabf;
sos_loop[0].somModel.sram_ptr[2][218]=2;
sos_loop[0].somModel.sram_dat[2][219][0]=96'hc8cd9;
sos_loop[0].somModel.sram_ptr[2][219]=2;
sos_loop[0].somModel.sram_dat[2][220][0]=96'h20926d;
sos_loop[0].somModel.sram_ptr[2][220]=2;
sos_loop[0].somModel.sram_dat[2][221][0]=96'hc358af;
sos_loop[0].somModel.sram_ptr[2][221]=2;
sos_loop[0].somModel.sram_dat[2][222][0]=96'h5bb9eb;
sos_loop[0].somModel.sram_ptr[2][222]=2;
sos_loop[0].somModel.sram_dat[2][223][0]=96'hb1e73e;
sos_loop[0].somModel.sram_ptr[2][223]=2;
sos_loop[0].somModel.sram_dat[2][224][0]=96'h591f46;
sos_loop[0].somModel.sram_ptr[2][224]=2;
sos_loop[0].somModel.sram_dat[2][225][0]=96'h7367d3;
sos_loop[0].somModel.sram_ptr[2][225]=2;
sos_loop[0].somModel.sram_dat[2][226][0]=96'h638b62;
sos_loop[0].somModel.sram_ptr[2][226]=2;
sos_loop[0].somModel.sram_dat[2][227][0]=96'h637b90;
sos_loop[0].somModel.sram_ptr[2][227]=2;
sos_loop[0].somModel.sram_dat[2][228][0]=96'h8d74b6;
sos_loop[0].somModel.sram_ptr[2][228]=2;
sos_loop[0].somModel.sram_dat[2][229][0]=96'h5c8f52;
sos_loop[0].somModel.sram_ptr[2][229]=2;
sos_loop[0].somModel.sram_dat[2][230][0]=96'hd7ee49;
sos_loop[0].somModel.sram_ptr[2][230]=2;
sos_loop[0].somModel.sram_dat[2][231][0]=96'hd72b91;
sos_loop[0].somModel.sram_ptr[2][231]=2;
sos_loop[0].somModel.sram_dat[2][232][0]=96'h816c24;
sos_loop[0].somModel.sram_ptr[2][232]=2;
sos_loop[0].somModel.sram_dat[2][233][0]=96'hde97a8;
sos_loop[0].somModel.sram_ptr[2][233]=2;
sos_loop[0].somModel.sram_dat[2][234][0]=96'h4ef26b;
sos_loop[0].somModel.sram_ptr[2][234]=2;
sos_loop[0].somModel.sram_dat[2][235][0]=96'hafbc7c;
sos_loop[0].somModel.sram_ptr[2][235]=2;
sos_loop[0].somModel.sram_dat[2][236][0]=96'h337d7d;
sos_loop[0].somModel.sram_ptr[2][236]=2;
sos_loop[0].somModel.sram_dat[2][237][0]=96'h781a2b;
sos_loop[0].somModel.sram_ptr[2][237]=2;
sos_loop[0].somModel.sram_dat[2][238][0]=96'hb4e99c;
sos_loop[0].somModel.sram_ptr[2][238]=2;
sos_loop[0].somModel.sram_dat[2][239][0]=96'ha1d931;
sos_loop[0].somModel.sram_ptr[2][239]=2;
sos_loop[0].somModel.sram_dat[2][240][0]=96'h2e3027;
sos_loop[0].somModel.sram_ptr[2][240]=2;
sos_loop[0].somModel.sram_dat[2][241][0]=96'hf983f9;
sos_loop[0].somModel.sram_ptr[2][241]=2;
sos_loop[0].somModel.sram_dat[2][242][0]=96'h56ed80;
sos_loop[0].somModel.sram_ptr[2][242]=2;
sos_loop[0].somModel.sram_dat[2][243][0]=96'h5200ab;
sos_loop[0].somModel.sram_ptr[2][243]=2;
sos_loop[0].somModel.sram_dat[2][244][0]=96'h637797;
sos_loop[0].somModel.sram_ptr[2][244]=2;
sos_loop[0].somModel.sram_dat[2][245][0]=96'hdd2137;
sos_loop[0].somModel.sram_ptr[2][245]=2;
sos_loop[0].somModel.sram_dat[2][246][0]=96'hfd2416;
sos_loop[0].somModel.sram_ptr[2][246]=2;
sos_loop[0].somModel.sram_dat[2][247][0]=96'hf3a4f0;
sos_loop[0].somModel.sram_ptr[2][247]=2;
sos_loop[0].somModel.sram_dat[2][248][0]=96'h44c886;
sos_loop[0].somModel.sram_ptr[2][248]=2;
sos_loop[0].somModel.sram_dat[2][249][0]=96'hceb410;
sos_loop[0].somModel.sram_ptr[2][249]=2;
sos_loop[0].somModel.sram_dat[2][250][0]=96'hf59b12;
sos_loop[0].somModel.sram_ptr[2][250]=2;
sos_loop[0].somModel.sram_dat[2][251][0]=96'he49bd0;
sos_loop[0].somModel.sram_ptr[2][251]=2;
sos_loop[0].somModel.sram_dat[2][252][0]=96'h638997;
sos_loop[0].somModel.sram_ptr[2][252]=2;
sos_loop[0].somModel.sram_dat[2][253][0]=96'h2f7580;
sos_loop[0].somModel.sram_ptr[2][253]=2;
sos_loop[0].somModel.sram_dat[2][254][0]=96'h1c10a8;
sos_loop[0].somModel.sram_ptr[2][254]=2;
sos_loop[0].somModel.sram_dat[2][255][0]=96'h879f04;
sos_loop[0].somModel.sram_ptr[2][255]=2;
sos_loop[0].somModel.sram_dat[2][256][0]=96'hbab2c4;
sos_loop[0].somModel.sram_ptr[2][256]=2;
sos_loop[0].somModel.sram_dat[2][257][0]=96'ha22715;
sos_loop[0].somModel.sram_ptr[2][257]=2;
sos_loop[0].somModel.sram_dat[2][258][0]=96'hf23b5e;
sos_loop[0].somModel.sram_ptr[2][258]=2;
sos_loop[0].somModel.sram_dat[2][259][0]=96'hfdc001;
sos_loop[0].somModel.sram_ptr[2][259]=2;
sos_loop[0].somModel.sram_dat[2][260][0]=96'h288bf0;
sos_loop[0].somModel.sram_ptr[2][260]=2;
sos_loop[0].somModel.sram_dat[2][261][0]=96'h662d40;
sos_loop[0].somModel.sram_ptr[2][261]=2;
sos_loop[0].somModel.sram_dat[2][262][0]=96'h72cef9;
sos_loop[0].somModel.sram_ptr[2][262]=2;
sos_loop[0].somModel.sram_dat[2][263][0]=96'h87666;
sos_loop[0].somModel.sram_ptr[2][263]=2;
sos_loop[0].somModel.sram_dat[2][264][0]=96'hf522c4;
sos_loop[0].somModel.sram_ptr[2][264]=2;
sos_loop[0].somModel.sram_dat[2][265][0]=96'hcf63c5;
sos_loop[0].somModel.sram_ptr[2][265]=2;
sos_loop[0].somModel.sram_dat[2][266][0]=96'he18e89;
sos_loop[0].somModel.sram_ptr[2][266]=2;
sos_loop[0].somModel.sram_dat[2][267][0]=96'ha2bc46;
sos_loop[0].somModel.sram_ptr[2][267]=2;
sos_loop[0].somModel.sram_dat[2][268][0]=96'h41996f;
sos_loop[0].somModel.sram_ptr[2][268]=2;
sos_loop[0].somModel.sram_dat[2][269][0]=96'h5e2a51;
sos_loop[0].somModel.sram_ptr[2][269]=2;
sos_loop[0].somModel.sram_dat[2][270][0]=96'h46b451;
sos_loop[0].somModel.sram_ptr[2][270]=2;
sos_loop[0].somModel.sram_dat[2][271][0]=96'hee2aae;
sos_loop[0].somModel.sram_ptr[2][271]=2;
sos_loop[0].somModel.sram_dat[2][272][0]=96'hb33948;
sos_loop[0].somModel.sram_ptr[2][272]=2;
sos_loop[0].somModel.sram_dat[2][273][0]=96'h7587fe;
sos_loop[0].somModel.sram_ptr[2][273]=2;
sos_loop[0].somModel.sram_dat[2][274][0]=96'h4584c5;
sos_loop[0].somModel.sram_ptr[2][274]=2;
sos_loop[0].somModel.sram_dat[2][275][0]=96'h4532c5;
sos_loop[0].somModel.sram_ptr[2][275]=2;
sos_loop[0].somModel.sram_dat[2][276][0]=96'h7754d8;
sos_loop[0].somModel.sram_ptr[2][276]=2;
sos_loop[0].somModel.sram_dat[2][277][0]=96'h2b77b;
sos_loop[0].somModel.sram_ptr[2][277]=2;
sos_loop[0].somModel.sram_dat[2][278][0]=96'h8f7473;
sos_loop[0].somModel.sram_ptr[2][278]=2;
sos_loop[0].somModel.sram_dat[2][279][0]=96'hff2471;
sos_loop[0].somModel.sram_ptr[2][279]=2;
sos_loop[0].somModel.sram_dat[2][280][0]=96'h14b05f;
sos_loop[0].somModel.sram_ptr[2][280]=2;
sos_loop[0].somModel.sram_dat[2][281][0]=96'hdf9570;
sos_loop[0].somModel.sram_ptr[2][281]=2;
sos_loop[0].somModel.sram_dat[2][282][0]=96'h153dbb;
sos_loop[0].somModel.sram_ptr[2][282]=2;
sos_loop[0].somModel.sram_dat[2][283][0]=96'hc5d62c;
sos_loop[0].somModel.sram_ptr[2][283]=2;
sos_loop[0].somModel.sram_dat[2][284][0]=96'h6bf1fb;
sos_loop[0].somModel.sram_ptr[2][284]=2;
sos_loop[0].somModel.sram_dat[2][285][0]=96'h25d7ea;
sos_loop[0].somModel.sram_ptr[2][285]=2;
sos_loop[0].somModel.sram_dat[2][286][0]=96'h7d1082;
sos_loop[0].somModel.sram_ptr[2][286]=2;
sos_loop[0].somModel.sram_dat[2][287][0]=96'h5f39c9;
sos_loop[0].somModel.sram_ptr[2][287]=2;
sos_loop[0].somModel.sram_dat[2][288][0]=96'h9fe99;
sos_loop[0].somModel.sram_ptr[2][288]=2;
sos_loop[0].somModel.sram_dat[2][289][0]=96'h7b04db;
sos_loop[0].somModel.sram_ptr[2][289]=2;
sos_loop[0].somModel.sram_dat[2][290][0]=96'h29dd6a;
sos_loop[0].somModel.sram_ptr[2][290]=2;
sos_loop[0].somModel.sram_dat[2][291][0]=96'h1fcd7e;
sos_loop[0].somModel.sram_ptr[2][291]=2;
sos_loop[0].somModel.sram_dat[2][292][0]=96'h5b635c;
sos_loop[0].somModel.sram_ptr[2][292]=2;
sos_loop[0].somModel.sram_dat[2][293][0]=96'h6eda0f;
sos_loop[0].somModel.sram_ptr[2][293]=2;
sos_loop[0].somModel.sram_dat[2][294][0]=96'hcef008;
sos_loop[0].somModel.sram_ptr[2][294]=2;
sos_loop[0].somModel.sram_dat[2][295][0]=96'h32dc5e;
sos_loop[0].somModel.sram_ptr[2][295]=2;
sos_loop[0].somModel.sram_dat[2][296][0]=96'h50586f;
sos_loop[0].somModel.sram_ptr[2][296]=2;
sos_loop[0].somModel.sram_dat[2][297][0]=96'h6dc367;
sos_loop[0].somModel.sram_ptr[2][297]=2;
sos_loop[0].somModel.sram_dat[2][298][0]=96'h9c1de1;
sos_loop[0].somModel.sram_ptr[2][298]=2;
sos_loop[0].somModel.sram_dat[2][299][0]=96'hfd77d3;
sos_loop[0].somModel.sram_ptr[2][299]=2;
sos_loop[0].somModel.sram_dat[2][300][0]=96'hd3c5d4;
sos_loop[0].somModel.sram_ptr[2][300]=2;
sos_loop[0].somModel.sram_dat[2][301][0]=96'hfdb0d;
sos_loop[0].somModel.sram_ptr[2][301]=2;
sos_loop[0].somModel.sram_dat[2][302][0]=96'h25d51;
sos_loop[0].somModel.sram_ptr[2][302]=2;
sos_loop[0].somModel.sram_dat[2][303][0]=96'he88800;
sos_loop[0].somModel.sram_ptr[2][303]=2;
sos_loop[0].somModel.sram_dat[2][304][0]=96'hc08b8e;
sos_loop[0].somModel.sram_ptr[2][304]=2;
sos_loop[0].somModel.sram_dat[2][305][0]=96'h3f0392;
sos_loop[0].somModel.sram_ptr[2][305]=2;
sos_loop[0].somModel.sram_dat[2][306][0]=96'ha02fb5;
sos_loop[0].somModel.sram_ptr[2][306]=2;
sos_loop[0].somModel.sram_dat[2][307][0]=96'h21607f;
sos_loop[0].somModel.sram_ptr[2][307]=2;
sos_loop[0].somModel.sram_dat[2][308][0]=96'h8f612f;
sos_loop[0].somModel.sram_ptr[2][308]=2;
sos_loop[0].somModel.sram_dat[2][309][0]=96'h34a36e;
sos_loop[0].somModel.sram_ptr[2][309]=2;
sos_loop[0].somModel.sram_dat[2][310][0]=96'h899446;
sos_loop[0].somModel.sram_ptr[2][310]=2;
sos_loop[0].somModel.sram_dat[2][311][0]=96'haeaee1;
sos_loop[0].somModel.sram_ptr[2][311]=2;
sos_loop[0].somModel.sram_dat[2][312][0]=96'hefa58;
sos_loop[0].somModel.sram_ptr[2][312]=2;
sos_loop[0].somModel.sram_dat[2][313][0]=96'h7c121d;
sos_loop[0].somModel.sram_ptr[2][313]=2;
sos_loop[0].somModel.sram_dat[2][314][0]=96'h84c243;
sos_loop[0].somModel.sram_ptr[2][314]=2;
sos_loop[0].somModel.sram_dat[2][315][0]=96'h6fa6f1;
sos_loop[0].somModel.sram_ptr[2][315]=2;
sos_loop[0].somModel.sram_dat[2][316][0]=96'he50d93;
sos_loop[0].somModel.sram_ptr[2][316]=2;
sos_loop[0].somModel.sram_dat[2][317][0]=96'h30a2f4;
sos_loop[0].somModel.sram_ptr[2][317]=2;
sos_loop[0].somModel.sram_dat[2][318][0]=96'h28773f;
sos_loop[0].somModel.sram_ptr[2][318]=2;
sos_loop[0].somModel.sram_dat[2][319][0]=96'h266b7;
sos_loop[0].somModel.sram_ptr[2][319]=2;
sos_loop[0].somModel.sram_dat[2][320][0]=96'ha9817d;
sos_loop[0].somModel.sram_ptr[2][320]=2;
sos_loop[0].somModel.sram_dat[2][321][0]=96'h3920db;
sos_loop[0].somModel.sram_ptr[2][321]=2;
sos_loop[0].somModel.sram_dat[2][322][0]=96'h3bfaad;
sos_loop[0].somModel.sram_ptr[2][322]=2;
sos_loop[0].somModel.sram_dat[2][323][0]=96'hd9c7f1;
sos_loop[0].somModel.sram_ptr[2][323]=2;
sos_loop[0].somModel.sram_dat[2][324][0]=96'h5c0486;
sos_loop[0].somModel.sram_ptr[2][324]=2;
sos_loop[0].somModel.sram_dat[2][325][0]=96'hd00200;
sos_loop[0].somModel.sram_ptr[2][325]=2;
sos_loop[0].somModel.sram_dat[2][326][0]=96'hd49869;
sos_loop[0].somModel.sram_ptr[2][326]=2;
sos_loop[0].somModel.sram_dat[2][327][0]=96'h89ee4e;
sos_loop[0].somModel.sram_ptr[2][327]=2;
sos_loop[0].somModel.sram_dat[2][328][0]=96'hdf942f;
sos_loop[0].somModel.sram_ptr[2][328]=2;
sos_loop[0].somModel.sram_dat[2][329][0]=96'h84601d;
sos_loop[0].somModel.sram_ptr[2][329]=2;
sos_loop[0].somModel.sram_dat[2][330][0]=96'h1808be;
sos_loop[0].somModel.sram_ptr[2][330]=2;
sos_loop[0].somModel.sram_dat[2][331][0]=96'hb502fb;
sos_loop[0].somModel.sram_ptr[2][331]=2;
sos_loop[0].somModel.sram_dat[2][332][0]=96'h9f2b20;
sos_loop[0].somModel.sram_ptr[2][332]=2;
sos_loop[0].somModel.sram_dat[2][333][0]=96'hb2fa64;
sos_loop[0].somModel.sram_ptr[2][333]=2;
sos_loop[0].somModel.sram_dat[2][334][0]=96'h80dd3b;
sos_loop[0].somModel.sram_ptr[2][334]=2;
sos_loop[0].somModel.sram_dat[2][335][0]=96'h38568a;
sos_loop[0].somModel.sram_ptr[2][335]=2;
sos_loop[0].somModel.sram_dat[2][336][0]=96'hea6666;
sos_loop[0].somModel.sram_ptr[2][336]=2;
sos_loop[0].somModel.sram_dat[2][337][0]=96'hdfa001;
sos_loop[0].somModel.sram_ptr[2][337]=2;
sos_loop[0].somModel.sram_dat[2][338][0]=96'h396ef;
sos_loop[0].somModel.sram_ptr[2][338]=2;
sos_loop[0].somModel.sram_dat[2][339][0]=96'h61ba43;
sos_loop[0].somModel.sram_ptr[2][339]=2;
sos_loop[0].somModel.sram_dat[2][340][0]=96'h80209;
sos_loop[0].somModel.sram_ptr[2][340]=2;
sos_loop[0].somModel.sram_dat[2][341][0]=96'h5b8fa1;
sos_loop[0].somModel.sram_ptr[2][341]=2;
sos_loop[0].somModel.sram_dat[2][342][0]=96'h61c5cc;
sos_loop[0].somModel.sram_ptr[2][342]=2;
sos_loop[0].somModel.sram_dat[2][343][0]=96'hb26ef1;
sos_loop[0].somModel.sram_ptr[2][343]=2;
sos_loop[0].somModel.sram_dat[2][344][0]=96'h407501;
sos_loop[0].somModel.sram_ptr[2][344]=2;
sos_loop[0].somModel.sram_dat[2][345][0]=96'h28ace5;
sos_loop[0].somModel.sram_ptr[2][345]=2;
sos_loop[0].somModel.sram_dat[2][346][0]=96'hc579b9;
sos_loop[0].somModel.sram_ptr[2][346]=2;
sos_loop[0].somModel.sram_dat[2][347][0]=96'h9bfb01;
sos_loop[0].somModel.sram_ptr[2][347]=2;
sos_loop[0].somModel.sram_dat[2][348][0]=96'hf34eb;
sos_loop[0].somModel.sram_ptr[2][348]=2;
sos_loop[0].somModel.sram_dat[2][349][0]=96'hab2f3d;
sos_loop[0].somModel.sram_ptr[2][349]=2;
sos_loop[0].somModel.sram_dat[2][350][0]=96'h186408;
sos_loop[0].somModel.sram_ptr[2][350]=2;
sos_loop[0].somModel.sram_dat[2][351][0]=96'h22a3c9;
sos_loop[0].somModel.sram_ptr[2][351]=2;
sos_loop[0].somModel.sram_dat[2][352][0]=96'h9aa041;
sos_loop[0].somModel.sram_ptr[2][352]=2;
sos_loop[0].somModel.sram_dat[2][353][0]=96'hb46f64;
sos_loop[0].somModel.sram_ptr[2][353]=2;
sos_loop[0].somModel.sram_dat[2][354][0]=96'h48548b;
sos_loop[0].somModel.sram_ptr[2][354]=2;
sos_loop[0].somModel.sram_dat[2][355][0]=96'he7ee30;
sos_loop[0].somModel.sram_ptr[2][355]=2;
sos_loop[0].somModel.sram_dat[2][356][0]=96'hc7e65;
sos_loop[0].somModel.sram_ptr[2][356]=2;
sos_loop[0].somModel.sram_dat[2][357][0]=96'hc4e05f;
sos_loop[0].somModel.sram_ptr[2][357]=2;
sos_loop[0].somModel.sram_dat[2][358][0]=96'hcdeb94;
sos_loop[0].somModel.sram_ptr[2][358]=2;
sos_loop[0].somModel.sram_dat[2][359][0]=96'hc6fbde;
sos_loop[0].somModel.sram_ptr[2][359]=2;
sos_loop[0].somModel.sram_dat[2][360][0]=96'h4364d2;
sos_loop[0].somModel.sram_ptr[2][360]=2;
sos_loop[0].somModel.sram_dat[2][361][0]=96'h54c878;
sos_loop[0].somModel.sram_ptr[2][361]=2;
sos_loop[0].somModel.sram_dat[2][362][0]=96'h244700;
sos_loop[0].somModel.sram_ptr[2][362]=2;
sos_loop[0].somModel.sram_dat[2][363][0]=96'h3a7f6d;
sos_loop[0].somModel.sram_ptr[2][363]=2;
sos_loop[0].somModel.sram_dat[2][364][0]=96'he03a58;
sos_loop[0].somModel.sram_ptr[2][364]=2;
sos_loop[0].somModel.sram_dat[2][365][0]=96'hb0efa4;
sos_loop[0].somModel.sram_ptr[2][365]=2;
sos_loop[0].somModel.sram_dat[2][366][0]=96'h1e6831;
sos_loop[0].somModel.sram_ptr[2][366]=2;
sos_loop[0].somModel.sram_dat[2][367][0]=96'h323acf;
sos_loop[0].somModel.sram_ptr[2][367]=2;
sos_loop[0].somModel.sram_dat[2][368][0]=96'h1ab23b;
sos_loop[0].somModel.sram_ptr[2][368]=2;
sos_loop[0].somModel.sram_dat[2][369][0]=96'h153918;
sos_loop[0].somModel.sram_ptr[2][369]=2;
sos_loop[0].somModel.sram_dat[2][370][0]=96'ha376d9;
sos_loop[0].somModel.sram_ptr[2][370]=2;
sos_loop[0].somModel.sram_dat[2][371][0]=96'h66c250;
sos_loop[0].somModel.sram_ptr[2][371]=2;
sos_loop[0].somModel.sram_dat[2][372][0]=96'hf46295;
sos_loop[0].somModel.sram_ptr[2][372]=2;
sos_loop[0].somModel.sram_dat[2][373][0]=96'h909a33;
sos_loop[0].somModel.sram_ptr[2][373]=2;
sos_loop[0].somModel.sram_dat[2][374][0]=96'hb903f6;
sos_loop[0].somModel.sram_ptr[2][374]=2;
sos_loop[0].somModel.sram_dat[2][375][0]=96'h876713;
sos_loop[0].somModel.sram_ptr[2][375]=2;
sos_loop[0].somModel.sram_dat[2][376][0]=96'hf203b1;
sos_loop[0].somModel.sram_ptr[2][376]=2;
sos_loop[0].somModel.sram_dat[2][377][0]=96'h7035e4;
sos_loop[0].somModel.sram_ptr[2][377]=2;
sos_loop[0].somModel.sram_dat[2][378][0]=96'he24033;
sos_loop[0].somModel.sram_ptr[2][378]=2;
sos_loop[0].somModel.sram_dat[2][379][0]=96'he8a4a2;
sos_loop[0].somModel.sram_ptr[2][379]=2;
sos_loop[0].somModel.sram_dat[2][380][0]=96'hece548;
sos_loop[0].somModel.sram_ptr[2][380]=2;
sos_loop[0].somModel.sram_dat[2][381][0]=96'h586dfc;
sos_loop[0].somModel.sram_ptr[2][381]=2;
sos_loop[0].somModel.sram_dat[2][382][0]=96'h8c1319;
sos_loop[0].somModel.sram_ptr[2][382]=2;
sos_loop[0].somModel.sram_dat[2][383][0]=96'h725176;
sos_loop[0].somModel.sram_ptr[2][383]=2;
sos_loop[0].somModel.sram_dat[2][384][0]=96'h56cec2;
sos_loop[0].somModel.sram_ptr[2][384]=2;
sos_loop[0].somModel.sram_dat[2][385][0]=96'h639a04;
sos_loop[0].somModel.sram_ptr[2][385]=2;
sos_loop[0].somModel.sram_dat[2][386][0]=96'h5327e0;
sos_loop[0].somModel.sram_ptr[2][386]=2;
sos_loop[0].somModel.sram_dat[2][387][0]=96'h1462c7;
sos_loop[0].somModel.sram_ptr[2][387]=2;
sos_loop[0].somModel.sram_dat[2][388][0]=96'hd89f5;
sos_loop[0].somModel.sram_ptr[2][388]=2;
sos_loop[0].somModel.sram_dat[2][389][0]=96'h3902ae;
sos_loop[0].somModel.sram_ptr[2][389]=2;
sos_loop[0].somModel.sram_dat[2][390][0]=96'ha2cbeb;
sos_loop[0].somModel.sram_ptr[2][390]=2;
sos_loop[0].somModel.sram_dat[2][391][0]=96'hf6681;
sos_loop[0].somModel.sram_ptr[2][391]=2;
sos_loop[0].somModel.sram_dat[2][392][0]=96'h5dcafd;
sos_loop[0].somModel.sram_ptr[2][392]=2;
sos_loop[0].somModel.sram_dat[2][393][0]=96'h691152;
sos_loop[0].somModel.sram_ptr[2][393]=2;
sos_loop[0].somModel.sram_dat[2][394][0]=96'h76bcf7;
sos_loop[0].somModel.sram_ptr[2][394]=2;
sos_loop[0].somModel.sram_dat[2][395][0]=96'h655333;
sos_loop[0].somModel.sram_ptr[2][395]=2;
sos_loop[0].somModel.sram_dat[2][396][0]=96'h67c107;
sos_loop[0].somModel.sram_ptr[2][396]=2;
sos_loop[0].somModel.sram_dat[2][397][0]=96'hbd651c;
sos_loop[0].somModel.sram_ptr[2][397]=2;
sos_loop[0].somModel.sram_dat[2][398][0]=96'hd88fbe;
sos_loop[0].somModel.sram_ptr[2][398]=2;
sos_loop[0].somModel.sram_dat[2][399][0]=96'h3fa26a;
sos_loop[0].somModel.sram_ptr[2][399]=2;
sos_loop[0].somModel.sram_dat[2][400][0]=96'hbe3762;
sos_loop[0].somModel.sram_ptr[2][400]=2;
sos_loop[0].somModel.sram_dat[2][401][0]=96'hee1fc4;
sos_loop[0].somModel.sram_ptr[2][401]=2;
sos_loop[0].somModel.sram_dat[2][402][0]=96'hb30bdf;
sos_loop[0].somModel.sram_ptr[2][402]=2;
sos_loop[0].somModel.sram_dat[2][403][0]=96'h977fec;
sos_loop[0].somModel.sram_ptr[2][403]=2;
sos_loop[0].somModel.sram_dat[2][404][0]=96'hf34eee;
sos_loop[0].somModel.sram_ptr[2][404]=2;
sos_loop[0].somModel.sram_dat[2][405][0]=96'h88c78e;
sos_loop[0].somModel.sram_ptr[2][405]=2;
sos_loop[0].somModel.sram_dat[2][406][0]=96'h50186a;
sos_loop[0].somModel.sram_ptr[2][406]=2;
sos_loop[0].somModel.sram_dat[2][407][0]=96'h22c496;
sos_loop[0].somModel.sram_ptr[2][407]=2;
sos_loop[0].somModel.sram_dat[2][408][0]=96'h74ba14;
sos_loop[0].somModel.sram_ptr[2][408]=2;
sos_loop[0].somModel.sram_dat[2][409][0]=96'h5fa922;
sos_loop[0].somModel.sram_ptr[2][409]=2;
sos_loop[0].somModel.sram_dat[2][410][0]=96'h9f94e;
sos_loop[0].somModel.sram_ptr[2][410]=2;
sos_loop[0].somModel.sram_dat[2][411][0]=96'h66d9fb;
sos_loop[0].somModel.sram_ptr[2][411]=2;
sos_loop[0].somModel.sram_dat[2][412][0]=96'h10bb50;
sos_loop[0].somModel.sram_ptr[2][412]=2;
sos_loop[0].somModel.sram_dat[2][413][0]=96'h139b8e;
sos_loop[0].somModel.sram_ptr[2][413]=2;
sos_loop[0].somModel.sram_dat[2][414][0]=96'h34094f;
sos_loop[0].somModel.sram_ptr[2][414]=2;
sos_loop[0].somModel.sram_dat[2][415][0]=96'hf852df;
sos_loop[0].somModel.sram_ptr[2][415]=2;
sos_loop[0].somModel.sram_dat[2][416][0]=96'hb4b4a5;
sos_loop[0].somModel.sram_ptr[2][416]=2;
sos_loop[0].somModel.sram_dat[2][417][0]=96'h7de478;
sos_loop[0].somModel.sram_ptr[2][417]=2;
sos_loop[0].somModel.sram_dat[2][418][0]=96'h3db18f;
sos_loop[0].somModel.sram_ptr[2][418]=2;
sos_loop[0].somModel.sram_dat[2][419][0]=96'hd272a2;
sos_loop[0].somModel.sram_ptr[2][419]=2;
sos_loop[0].somModel.sram_dat[2][420][0]=96'h8fb4b5;
sos_loop[0].somModel.sram_ptr[2][420]=2;
sos_loop[0].somModel.sram_dat[2][421][0]=96'h39e1a2;
sos_loop[0].somModel.sram_ptr[2][421]=2;
sos_loop[0].somModel.sram_dat[2][422][0]=96'hbcc07b;
sos_loop[0].somModel.sram_ptr[2][422]=2;
sos_loop[0].somModel.sram_dat[2][423][0]=96'hb2ab05;
sos_loop[0].somModel.sram_ptr[2][423]=2;
sos_loop[0].somModel.sram_dat[2][424][0]=96'hf3b478;
sos_loop[0].somModel.sram_ptr[2][424]=2;
sos_loop[0].somModel.sram_dat[2][425][0]=96'h9c9331;
sos_loop[0].somModel.sram_ptr[2][425]=2;
sos_loop[0].somModel.sram_dat[2][426][0]=96'h570f8;
sos_loop[0].somModel.sram_ptr[2][426]=2;
sos_loop[0].somModel.sram_dat[2][427][0]=96'h92489c;
sos_loop[0].somModel.sram_ptr[2][427]=2;
sos_loop[0].somModel.sram_dat[2][428][0]=96'hd0fc4d;
sos_loop[0].somModel.sram_ptr[2][428]=2;
sos_loop[0].somModel.sram_dat[2][429][0]=96'h2acd7b;
sos_loop[0].somModel.sram_ptr[2][429]=2;
sos_loop[0].somModel.sram_dat[2][430][0]=96'hab42dd;
sos_loop[0].somModel.sram_ptr[2][430]=2;
sos_loop[0].somModel.sram_dat[2][431][0]=96'he77e1b;
sos_loop[0].somModel.sram_ptr[2][431]=2;
sos_loop[0].somModel.sram_dat[2][432][0]=96'h81a3c5;
sos_loop[0].somModel.sram_ptr[2][432]=2;
sos_loop[0].somModel.sram_dat[2][433][0]=96'h6cf1fa;
sos_loop[0].somModel.sram_ptr[2][433]=2;
sos_loop[0].somModel.sram_dat[2][434][0]=96'h34d05e;
sos_loop[0].somModel.sram_ptr[2][434]=2;
sos_loop[0].somModel.sram_dat[2][435][0]=96'h2b443d;
sos_loop[0].somModel.sram_ptr[2][435]=2;
sos_loop[0].somModel.sram_dat[2][436][0]=96'h97d73f;
sos_loop[0].somModel.sram_ptr[2][436]=2;
sos_loop[0].somModel.sram_dat[2][437][0]=96'h158478;
sos_loop[0].somModel.sram_ptr[2][437]=2;
sos_loop[0].somModel.sram_dat[2][438][0]=96'he145aa;
sos_loop[0].somModel.sram_ptr[2][438]=2;
sos_loop[0].somModel.sram_dat[2][439][0]=96'h1c385e;
sos_loop[0].somModel.sram_ptr[2][439]=2;
sos_loop[0].somModel.sram_dat[2][440][0]=96'hadbce3;
sos_loop[0].somModel.sram_ptr[2][440]=2;
sos_loop[0].somModel.sram_dat[2][441][0]=96'hd72c20;
sos_loop[0].somModel.sram_ptr[2][441]=2;
sos_loop[0].somModel.sram_dat[2][442][0]=96'h5a3b1b;
sos_loop[0].somModel.sram_ptr[2][442]=2;
sos_loop[0].somModel.sram_dat[2][443][0]=96'h5eaede;
sos_loop[0].somModel.sram_ptr[2][443]=2;
sos_loop[0].somModel.sram_dat[2][444][0]=96'h651848;
sos_loop[0].somModel.sram_ptr[2][444]=2;
sos_loop[0].somModel.sram_dat[2][445][0]=96'h977b39;
sos_loop[0].somModel.sram_ptr[2][445]=2;
sos_loop[0].somModel.sram_dat[2][446][0]=96'h5cea8e;
sos_loop[0].somModel.sram_ptr[2][446]=2;
sos_loop[0].somModel.sram_dat[2][447][0]=96'h3b6c9a;
sos_loop[0].somModel.sram_ptr[2][447]=2;
sos_loop[0].somModel.sram_dat[2][448][0]=96'h492ee4;
sos_loop[0].somModel.sram_ptr[2][448]=2;
sos_loop[0].somModel.sram_dat[2][449][0]=96'h9a047c;
sos_loop[0].somModel.sram_ptr[2][449]=2;
sos_loop[0].somModel.sram_dat[2][450][0]=96'h608036;
sos_loop[0].somModel.sram_ptr[2][450]=2;
sos_loop[0].somModel.sram_dat[2][451][0]=96'hcbe70e;
sos_loop[0].somModel.sram_ptr[2][451]=2;
sos_loop[0].somModel.sram_dat[2][452][0]=96'h1eb27a;
sos_loop[0].somModel.sram_ptr[2][452]=2;
sos_loop[0].somModel.sram_dat[2][453][0]=96'h751c3a;
sos_loop[0].somModel.sram_ptr[2][453]=2;
sos_loop[0].somModel.sram_dat[2][454][0]=96'h2b749f;
sos_loop[0].somModel.sram_ptr[2][454]=2;
sos_loop[0].somModel.sram_dat[2][455][0]=96'h7ab9cd;
sos_loop[0].somModel.sram_ptr[2][455]=2;
sos_loop[0].somModel.sram_dat[2][456][0]=96'hdb74b0;
sos_loop[0].somModel.sram_ptr[2][456]=2;
sos_loop[0].somModel.sram_dat[2][457][0]=96'h38ccf5;
sos_loop[0].somModel.sram_ptr[2][457]=2;
sos_loop[0].somModel.sram_dat[2][458][0]=96'hb81901;
sos_loop[0].somModel.sram_ptr[2][458]=2;
sos_loop[0].somModel.sram_dat[2][459][0]=96'hdb6f8a;
sos_loop[0].somModel.sram_ptr[2][459]=2;
sos_loop[0].somModel.sram_dat[2][460][0]=96'hbdfaee;
sos_loop[0].somModel.sram_ptr[2][460]=2;
sos_loop[0].somModel.sram_dat[2][461][0]=96'hab9134;
sos_loop[0].somModel.sram_ptr[2][461]=2;
sos_loop[0].somModel.sram_dat[2][462][0]=96'h6d74aa;
sos_loop[0].somModel.sram_ptr[2][462]=2;
sos_loop[0].somModel.sram_dat[2][463][0]=96'hf71076;
sos_loop[0].somModel.sram_ptr[2][463]=2;
sos_loop[0].somModel.sram_dat[2][464][0]=96'h579bdc;
sos_loop[0].somModel.sram_ptr[2][464]=2;
sos_loop[0].somModel.sram_dat[2][465][0]=96'hbbbd64;
sos_loop[0].somModel.sram_ptr[2][465]=2;
sos_loop[0].somModel.sram_dat[2][466][0]=96'h83ae74;
sos_loop[0].somModel.sram_ptr[2][466]=2;
sos_loop[0].somModel.sram_dat[2][467][0]=96'hf8c1d9;
sos_loop[0].somModel.sram_ptr[2][467]=2;
sos_loop[0].somModel.sram_dat[2][468][0]=96'hc8ed3e;
sos_loop[0].somModel.sram_ptr[2][468]=2;
sos_loop[0].somModel.sram_dat[2][469][0]=96'h2bf8dc;
sos_loop[0].somModel.sram_ptr[2][469]=2;
sos_loop[0].somModel.sram_dat[2][470][0]=96'h16e5de;
sos_loop[0].somModel.sram_ptr[2][470]=2;
sos_loop[0].somModel.sram_dat[2][471][0]=96'hb99492;
sos_loop[0].somModel.sram_ptr[2][471]=2;
sos_loop[0].somModel.sram_dat[2][472][0]=96'h820b16;
sos_loop[0].somModel.sram_ptr[2][472]=2;
sos_loop[0].somModel.sram_dat[2][473][0]=96'h8ae9cf;
sos_loop[0].somModel.sram_ptr[2][473]=2;
sos_loop[0].somModel.sram_dat[2][474][0]=96'hf6aad1;
sos_loop[0].somModel.sram_ptr[2][474]=2;
sos_loop[0].somModel.sram_dat[2][475][0]=96'hdef433;
sos_loop[0].somModel.sram_ptr[2][475]=2;
sos_loop[0].somModel.sram_dat[2][476][0]=96'h60e02b;
sos_loop[0].somModel.sram_ptr[2][476]=2;
sos_loop[0].somModel.sram_dat[2][477][0]=96'hba10d9;
sos_loop[0].somModel.sram_ptr[2][477]=2;
sos_loop[0].somModel.sram_dat[2][478][0]=96'h125ae0;
sos_loop[0].somModel.sram_ptr[2][478]=2;
sos_loop[0].somModel.sram_dat[2][479][0]=96'h75abca;
sos_loop[0].somModel.sram_ptr[2][479]=2;
sos_loop[0].somModel.sram_dat[2][480][0]=96'h7d0a37;
sos_loop[0].somModel.sram_ptr[2][480]=2;
sos_loop[0].somModel.sram_dat[2][481][0]=96'h76c3eb;
sos_loop[0].somModel.sram_ptr[2][481]=2;
sos_loop[0].somModel.sram_dat[2][482][0]=96'hee5867;
sos_loop[0].somModel.sram_ptr[2][482]=2;
sos_loop[0].somModel.sram_dat[2][483][0]=96'ha63aa9;
sos_loop[0].somModel.sram_ptr[2][483]=2;
sos_loop[0].somModel.sram_dat[2][484][0]=96'h3bf1a7;
sos_loop[0].somModel.sram_ptr[2][484]=2;
sos_loop[0].somModel.sram_dat[2][485][0]=96'h41b00e;
sos_loop[0].somModel.sram_ptr[2][485]=2;
sos_loop[0].somModel.sram_dat[2][486][0]=96'h5dfcea;
sos_loop[0].somModel.sram_ptr[2][486]=2;
sos_loop[0].somModel.sram_dat[2][487][0]=96'h856939;
sos_loop[0].somModel.sram_ptr[2][487]=2;
sos_loop[0].somModel.sram_dat[2][488][0]=96'h7fdd0;
sos_loop[0].somModel.sram_ptr[2][488]=2;
sos_loop[0].somModel.sram_dat[2][489][0]=96'hcac855;
sos_loop[0].somModel.sram_ptr[2][489]=2;
sos_loop[0].somModel.sram_dat[2][490][0]=96'h82c86b;
sos_loop[0].somModel.sram_ptr[2][490]=2;
sos_loop[0].somModel.sram_dat[2][491][0]=96'h7d64e0;
sos_loop[0].somModel.sram_ptr[2][491]=2;
sos_loop[0].somModel.sram_dat[2][492][0]=96'hc05790;
sos_loop[0].somModel.sram_ptr[2][492]=2;
sos_loop[0].somModel.sram_dat[2][493][0]=96'h41b488;
sos_loop[0].somModel.sram_ptr[2][493]=2;
sos_loop[0].somModel.sram_dat[2][494][0]=96'h19ef12;
sos_loop[0].somModel.sram_ptr[2][494]=2;
sos_loop[0].somModel.sram_dat[2][495][0]=96'h89d14b;
sos_loop[0].somModel.sram_ptr[2][495]=2;
sos_loop[0].somModel.sram_dat[2][496][0]=96'hb42732;
sos_loop[0].somModel.sram_ptr[2][496]=2;
sos_loop[0].somModel.sram_dat[2][497][0]=96'ha795fa;
sos_loop[0].somModel.sram_ptr[2][497]=2;
sos_loop[0].somModel.sram_dat[2][498][0]=96'ha72e70;
sos_loop[0].somModel.sram_ptr[2][498]=2;
sos_loop[0].somModel.sram_dat[2][499][0]=96'ha16e73;
sos_loop[0].somModel.sram_ptr[2][499]=2;
sos_loop[0].somModel.sram_dat[2][500][0]=96'h80fe5c;
sos_loop[0].somModel.sram_ptr[2][500]=2;
sos_loop[0].somModel.sram_dat[2][501][0]=96'hbdf1f7;
sos_loop[0].somModel.sram_ptr[2][501]=2;
sos_loop[0].somModel.sram_dat[2][502][0]=96'h24e03d;
sos_loop[0].somModel.sram_ptr[2][502]=2;
sos_loop[0].somModel.sram_dat[2][503][0]=96'hcd8833;
sos_loop[0].somModel.sram_ptr[2][503]=2;
sos_loop[0].somModel.sram_dat[2][504][0]=96'hd48427;
sos_loop[0].somModel.sram_ptr[2][504]=2;
sos_loop[0].somModel.sram_dat[2][505][0]=96'h29413e;
sos_loop[0].somModel.sram_ptr[2][505]=2;
sos_loop[0].somModel.sram_dat[2][506][0]=96'h99f215;
sos_loop[0].somModel.sram_ptr[2][506]=2;
sos_loop[0].somModel.sram_dat[2][507][0]=96'h43ea2c;
sos_loop[0].somModel.sram_ptr[2][507]=2;
sos_loop[0].somModel.sram_dat[2][508][0]=96'hb05ed6;
sos_loop[0].somModel.sram_ptr[2][508]=2;
sos_loop[0].somModel.sram_dat[2][509][0]=96'h359c4e;
sos_loop[0].somModel.sram_ptr[2][509]=2;
sos_loop[0].somModel.sram_dat[2][510][0]=96'ha53a50;
sos_loop[0].somModel.sram_ptr[2][510]=2;
sos_loop[0].somModel.sram_dat[2][511][0]=96'hba0217;
sos_loop[0].somModel.sram_ptr[2][511]=2;
sos_loop[0].somModel.sram_dat[2][512][0]=96'ha7a8be;
sos_loop[0].somModel.sram_ptr[2][512]=2;
sos_loop[0].somModel.sram_dat[2][513][0]=96'h117261;
sos_loop[0].somModel.sram_ptr[2][513]=2;
sos_loop[0].somModel.sram_dat[2][514][0]=96'hba40b1;
sos_loop[0].somModel.sram_ptr[2][514]=2;
sos_loop[0].somModel.sram_dat[2][515][0]=96'hd3778c;
sos_loop[0].somModel.sram_ptr[2][515]=2;
sos_loop[0].somModel.sram_dat[2][516][0]=96'h133300;
sos_loop[0].somModel.sram_ptr[2][516]=2;
sos_loop[0].somModel.sram_dat[2][517][0]=96'h8026d0;
sos_loop[0].somModel.sram_ptr[2][517]=2;
sos_loop[0].somModel.sram_dat[2][518][0]=96'h3c2a96;
sos_loop[0].somModel.sram_ptr[2][518]=2;
sos_loop[0].somModel.sram_dat[2][519][0]=96'haf2172;
sos_loop[0].somModel.sram_ptr[2][519]=2;
sos_loop[0].somModel.sram_dat[2][520][0]=96'hf83e69;
sos_loop[0].somModel.sram_ptr[2][520]=2;
sos_loop[0].somModel.sram_dat[2][521][0]=96'h2bae72;
sos_loop[0].somModel.sram_ptr[2][521]=2;
sos_loop[0].somModel.sram_dat[2][522][0]=96'haaffe3;
sos_loop[0].somModel.sram_ptr[2][522]=2;
sos_loop[0].somModel.sram_dat[2][523][0]=96'he47a3a;
sos_loop[0].somModel.sram_ptr[2][523]=2;
sos_loop[0].somModel.sram_dat[2][524][0]=96'hecf185;
sos_loop[0].somModel.sram_ptr[2][524]=2;
sos_loop[0].somModel.sram_dat[2][525][0]=96'h2ed0f5;
sos_loop[0].somModel.sram_ptr[2][525]=2;
sos_loop[0].somModel.sram_dat[2][526][0]=96'hd53425;
sos_loop[0].somModel.sram_ptr[2][526]=2;
sos_loop[0].somModel.sram_dat[2][527][0]=96'hecfd2a;
sos_loop[0].somModel.sram_ptr[2][527]=2;
sos_loop[0].somModel.sram_dat[2][528][0]=96'hc133a2;
sos_loop[0].somModel.sram_ptr[2][528]=2;
sos_loop[0].somModel.sram_dat[2][529][0]=96'hb51947;
sos_loop[0].somModel.sram_ptr[2][529]=2;
sos_loop[0].somModel.sram_dat[2][530][0]=96'h1f5b10;
sos_loop[0].somModel.sram_ptr[2][530]=2;
sos_loop[0].somModel.sram_dat[2][531][0]=96'h724175;
sos_loop[0].somModel.sram_ptr[2][531]=2;
sos_loop[0].somModel.sram_dat[2][532][0]=96'h4a6946;
sos_loop[0].somModel.sram_ptr[2][532]=2;
sos_loop[0].somModel.sram_dat[2][533][0]=96'hf4634a;
sos_loop[0].somModel.sram_ptr[2][533]=2;
sos_loop[0].somModel.sram_dat[2][534][0]=96'h74e5f6;
sos_loop[0].somModel.sram_ptr[2][534]=2;
sos_loop[0].somModel.sram_dat[2][535][0]=96'hb53980;
sos_loop[0].somModel.sram_ptr[2][535]=2;
sos_loop[0].somModel.sram_dat[2][536][0]=96'hbbd32a;
sos_loop[0].somModel.sram_ptr[2][536]=2;
sos_loop[0].somModel.sram_dat[2][537][0]=96'h4beff2;
sos_loop[0].somModel.sram_ptr[2][537]=2;
sos_loop[0].somModel.sram_dat[2][538][0]=96'hc8358f;
sos_loop[0].somModel.sram_ptr[2][538]=2;
sos_loop[0].somModel.sram_dat[2][539][0]=96'hcb9cd4;
sos_loop[0].somModel.sram_ptr[2][539]=2;
sos_loop[0].somModel.sram_dat[2][540][0]=96'h5a3371;
sos_loop[0].somModel.sram_ptr[2][540]=2;
sos_loop[0].somModel.sram_dat[2][541][0]=96'hb24300;
sos_loop[0].somModel.sram_ptr[2][541]=2;
sos_loop[0].somModel.sram_dat[2][542][0]=96'h1fb996;
sos_loop[0].somModel.sram_ptr[2][542]=2;
sos_loop[0].somModel.sram_dat[2][543][0]=96'hbd4f61;
sos_loop[0].somModel.sram_ptr[2][543]=2;
sos_loop[0].somModel.sram_dat[2][544][0]=96'h8abbcd;
sos_loop[0].somModel.sram_ptr[2][544]=2;
sos_loop[0].somModel.sram_dat[2][545][0]=96'hb9b2c6;
sos_loop[0].somModel.sram_ptr[2][545]=2;
sos_loop[0].somModel.sram_dat[2][546][0]=96'h638408;
sos_loop[0].somModel.sram_ptr[2][546]=2;
sos_loop[0].somModel.sram_dat[2][547][0]=96'hd821e0;
sos_loop[0].somModel.sram_ptr[2][547]=2;
sos_loop[0].somModel.sram_dat[2][548][0]=96'h694d89;
sos_loop[0].somModel.sram_ptr[2][548]=2;
sos_loop[0].somModel.sram_dat[2][549][0]=96'hcc2430;
sos_loop[0].somModel.sram_ptr[2][549]=2;
sos_loop[0].somModel.sram_dat[2][550][0]=96'hb3c95;
sos_loop[0].somModel.sram_ptr[2][550]=2;
sos_loop[0].somModel.sram_dat[2][551][0]=96'h2c40c9;
sos_loop[0].somModel.sram_ptr[2][551]=2;
sos_loop[0].somModel.sram_dat[2][552][0]=96'hec7053;
sos_loop[0].somModel.sram_ptr[2][552]=2;
sos_loop[0].somModel.sram_dat[2][553][0]=96'h8adfbd;
sos_loop[0].somModel.sram_ptr[2][553]=2;
sos_loop[0].somModel.sram_dat[2][554][0]=96'h15e421;
sos_loop[0].somModel.sram_ptr[2][554]=2;
sos_loop[0].somModel.sram_dat[2][555][0]=96'hcd639d;
sos_loop[0].somModel.sram_ptr[2][555]=2;
sos_loop[0].somModel.sram_dat[2][556][0]=96'h6a5ec;
sos_loop[0].somModel.sram_ptr[2][556]=2;
sos_loop[0].somModel.sram_dat[2][557][0]=96'h4837b3;
sos_loop[0].somModel.sram_ptr[2][557]=2;
sos_loop[0].somModel.sram_dat[2][558][0]=96'h3c1296;
sos_loop[0].somModel.sram_ptr[2][558]=2;
sos_loop[0].somModel.sram_dat[2][559][0]=96'h9854db;
sos_loop[0].somModel.sram_ptr[2][559]=2;
sos_loop[0].somModel.sram_dat[2][560][0]=96'he23953;
sos_loop[0].somModel.sram_ptr[2][560]=2;
sos_loop[0].somModel.sram_dat[2][561][0]=96'h6e5f61;
sos_loop[0].somModel.sram_ptr[2][561]=2;
sos_loop[0].somModel.sram_dat[2][562][0]=96'hb67704;
sos_loop[0].somModel.sram_ptr[2][562]=2;
sos_loop[0].somModel.sram_dat[2][563][0]=96'hc188f5;
sos_loop[0].somModel.sram_ptr[2][563]=2;
sos_loop[0].somModel.sram_dat[2][564][0]=96'h9f0af0;
sos_loop[0].somModel.sram_ptr[2][564]=2;
sos_loop[0].somModel.sram_dat[2][565][0]=96'h13deba;
sos_loop[0].somModel.sram_ptr[2][565]=2;
sos_loop[0].somModel.sram_dat[2][566][0]=96'hd836a2;
sos_loop[0].somModel.sram_ptr[2][566]=2;
sos_loop[0].somModel.sram_dat[2][567][0]=96'h378015;
sos_loop[0].somModel.sram_ptr[2][567]=2;
sos_loop[0].somModel.sram_dat[2][568][0]=96'h6857c;
sos_loop[0].somModel.sram_ptr[2][568]=2;
sos_loop[0].somModel.sram_dat[2][569][0]=96'h920848;
sos_loop[0].somModel.sram_ptr[2][569]=2;
sos_loop[0].somModel.sram_dat[2][570][0]=96'hdf91e5;
sos_loop[0].somModel.sram_ptr[2][570]=2;
sos_loop[0].somModel.sram_dat[2][571][0]=96'h203539;
sos_loop[0].somModel.sram_ptr[2][571]=2;
sos_loop[0].somModel.sram_dat[2][572][0]=96'he0e16e;
sos_loop[0].somModel.sram_ptr[2][572]=2;
sos_loop[0].somModel.sram_dat[2][573][0]=96'h518348;
sos_loop[0].somModel.sram_ptr[2][573]=2;
sos_loop[0].somModel.sram_dat[2][574][0]=96'h29589f;
sos_loop[0].somModel.sram_ptr[2][574]=2;
sos_loop[0].somModel.sram_dat[2][575][0]=96'hd5eff5;
sos_loop[0].somModel.sram_ptr[2][575]=2;
sos_loop[0].somModel.sram_dat[2][576][0]=96'ha8909a;
sos_loop[0].somModel.sram_ptr[2][576]=2;
sos_loop[0].somModel.sram_dat[2][577][0]=96'hc6ccb7;
sos_loop[0].somModel.sram_ptr[2][577]=2;
sos_loop[0].somModel.sram_dat[2][578][0]=96'h8fd56d;
sos_loop[0].somModel.sram_ptr[2][578]=2;
sos_loop[0].somModel.sram_dat[2][579][0]=96'hbf7f6d;
sos_loop[0].somModel.sram_ptr[2][579]=2;
sos_loop[0].somModel.sram_dat[2][580][0]=96'h6a229b;
sos_loop[0].somModel.sram_ptr[2][580]=2;
sos_loop[0].somModel.sram_dat[2][581][0]=96'ha7dd84;
sos_loop[0].somModel.sram_ptr[2][581]=2;
sos_loop[0].somModel.sram_dat[2][582][0]=96'h3d9854;
sos_loop[0].somModel.sram_ptr[2][582]=2;
sos_loop[0].somModel.sram_dat[2][583][0]=96'h3c87c6;
sos_loop[0].somModel.sram_ptr[2][583]=2;
sos_loop[0].somModel.sram_dat[2][584][0]=96'h588ad5;
sos_loop[0].somModel.sram_ptr[2][584]=2;
sos_loop[0].somModel.sram_dat[2][585][0]=96'heaaf14;
sos_loop[0].somModel.sram_ptr[2][585]=2;
sos_loop[0].somModel.sram_dat[2][586][0]=96'h344bf2;
sos_loop[0].somModel.sram_ptr[2][586]=2;
sos_loop[0].somModel.sram_dat[2][587][0]=96'h3d9161;
sos_loop[0].somModel.sram_ptr[2][587]=2;
sos_loop[0].somModel.sram_dat[2][588][0]=96'h415ce;
sos_loop[0].somModel.sram_ptr[2][588]=2;
sos_loop[0].somModel.sram_dat[2][589][0]=96'hb69cc;
sos_loop[0].somModel.sram_ptr[2][589]=2;
sos_loop[0].somModel.sram_dat[2][590][0]=96'hfe9312;
sos_loop[0].somModel.sram_ptr[2][590]=2;
sos_loop[0].somModel.sram_dat[2][591][0]=96'h878cb6;
sos_loop[0].somModel.sram_ptr[2][591]=2;
sos_loop[0].somModel.sram_dat[2][592][0]=96'h38cf4e;
sos_loop[0].somModel.sram_ptr[2][592]=2;
sos_loop[0].somModel.sram_dat[2][593][0]=96'h76dcb4;
sos_loop[0].somModel.sram_ptr[2][593]=2;
sos_loop[0].somModel.sram_dat[2][594][0]=96'h702f85;
sos_loop[0].somModel.sram_ptr[2][594]=2;
sos_loop[0].somModel.sram_dat[2][595][0]=96'hecdc20;
sos_loop[0].somModel.sram_ptr[2][595]=2;
sos_loop[0].somModel.sram_dat[2][596][0]=96'h64eed;
sos_loop[0].somModel.sram_ptr[2][596]=2;
sos_loop[0].somModel.sram_dat[2][597][0]=96'h197ad7;
sos_loop[0].somModel.sram_ptr[2][597]=2;
sos_loop[0].somModel.sram_dat[2][598][0]=96'h860fe2;
sos_loop[0].somModel.sram_ptr[2][598]=2;
sos_loop[0].somModel.sram_dat[2][599][0]=96'haafcfa;
sos_loop[0].somModel.sram_ptr[2][599]=2;
sos_loop[0].somModel.sram_dat[2][600][0]=96'hb3fdf0;
sos_loop[0].somModel.sram_ptr[2][600]=2;
sos_loop[0].somModel.sram_dat[2][601][0]=96'h75513;
sos_loop[0].somModel.sram_ptr[2][601]=2;
sos_loop[0].somModel.sram_dat[2][602][0]=96'h13141b;
sos_loop[0].somModel.sram_ptr[2][602]=2;
sos_loop[0].somModel.sram_dat[2][603][0]=96'hd07c80;
sos_loop[0].somModel.sram_ptr[2][603]=2;
sos_loop[0].somModel.sram_dat[2][604][0]=96'h7023d5;
sos_loop[0].somModel.sram_ptr[2][604]=2;
sos_loop[0].somModel.sram_dat[2][605][0]=96'h88bbc7;
sos_loop[0].somModel.sram_ptr[2][605]=2;
sos_loop[0].somModel.sram_dat[2][606][0]=96'h8bd1c2;
sos_loop[0].somModel.sram_ptr[2][606]=2;
sos_loop[0].somModel.sram_dat[2][607][0]=96'hede0cc;
sos_loop[0].somModel.sram_ptr[2][607]=2;
sos_loop[0].somModel.sram_dat[2][608][0]=96'h11d1b8;
sos_loop[0].somModel.sram_ptr[2][608]=2;
sos_loop[0].somModel.sram_dat[2][609][0]=96'hd0feb3;
sos_loop[0].somModel.sram_ptr[2][609]=2;
sos_loop[0].somModel.sram_dat[2][610][0]=96'hef7aab;
sos_loop[0].somModel.sram_ptr[2][610]=2;
sos_loop[0].somModel.sram_dat[2][611][0]=96'h929846;
sos_loop[0].somModel.sram_ptr[2][611]=2;
sos_loop[0].somModel.sram_dat[2][612][0]=96'h87f8f5;
sos_loop[0].somModel.sram_ptr[2][612]=2;
sos_loop[0].somModel.sram_dat[2][613][0]=96'hf6d906;
sos_loop[0].somModel.sram_ptr[2][613]=2;
sos_loop[0].somModel.sram_dat[2][614][0]=96'h301023;
sos_loop[0].somModel.sram_ptr[2][614]=2;
sos_loop[0].somModel.sram_dat[2][615][0]=96'hc0367e;
sos_loop[0].somModel.sram_ptr[2][615]=2;
sos_loop[0].somModel.sram_dat[2][616][0]=96'hb5225;
sos_loop[0].somModel.sram_ptr[2][616]=2;
sos_loop[0].somModel.sram_dat[2][617][0]=96'h1abda8;
sos_loop[0].somModel.sram_ptr[2][617]=2;
sos_loop[0].somModel.sram_dat[2][618][0]=96'hf76cf7;
sos_loop[0].somModel.sram_ptr[2][618]=2;
sos_loop[0].somModel.sram_dat[2][619][0]=96'h715672;
sos_loop[0].somModel.sram_ptr[2][619]=2;
sos_loop[0].somModel.sram_dat[2][620][0]=96'h7a6132;
sos_loop[0].somModel.sram_ptr[2][620]=2;
sos_loop[0].somModel.sram_dat[2][621][0]=96'h443d93;
sos_loop[0].somModel.sram_ptr[2][621]=2;
sos_loop[0].somModel.sram_dat[2][622][0]=96'heb213b;
sos_loop[0].somModel.sram_ptr[2][622]=2;
sos_loop[0].somModel.sram_dat[2][623][0]=96'h4d47a0;
sos_loop[0].somModel.sram_ptr[2][623]=2;
sos_loop[0].somModel.sram_dat[2][624][0]=96'ha05377;
sos_loop[0].somModel.sram_ptr[2][624]=2;
sos_loop[0].somModel.sram_dat[2][625][0]=96'h6ac1b8;
sos_loop[0].somModel.sram_ptr[2][625]=2;
sos_loop[0].somModel.sram_dat[2][626][0]=96'h7a773d;
sos_loop[0].somModel.sram_ptr[2][626]=2;
sos_loop[0].somModel.sram_dat[2][627][0]=96'he5e3a5;
sos_loop[0].somModel.sram_ptr[2][627]=2;
sos_loop[0].somModel.sram_dat[2][628][0]=96'hc9746b;
sos_loop[0].somModel.sram_ptr[2][628]=2;
sos_loop[0].somModel.sram_dat[2][629][0]=96'h23a9d3;
sos_loop[0].somModel.sram_ptr[2][629]=2;
sos_loop[0].somModel.sram_dat[2][630][0]=96'h4ec356;
sos_loop[0].somModel.sram_ptr[2][630]=2;
sos_loop[0].somModel.sram_dat[2][631][0]=96'h75d68;
sos_loop[0].somModel.sram_ptr[2][631]=2;
sos_loop[0].somModel.sram_dat[2][632][0]=96'h3f8eba;
sos_loop[0].somModel.sram_ptr[2][632]=2;
sos_loop[0].somModel.sram_dat[2][633][0]=96'h4d98e8;
sos_loop[0].somModel.sram_ptr[2][633]=2;
sos_loop[0].somModel.sram_dat[2][634][0]=96'h98da92;
sos_loop[0].somModel.sram_ptr[2][634]=2;
sos_loop[0].somModel.sram_dat[2][635][0]=96'hca02ef;
sos_loop[0].somModel.sram_ptr[2][635]=2;
sos_loop[0].somModel.sram_dat[2][636][0]=96'h924656;
sos_loop[0].somModel.sram_ptr[2][636]=2;
sos_loop[0].somModel.sram_dat[2][637][0]=96'h4eb306;
sos_loop[0].somModel.sram_ptr[2][637]=2;
sos_loop[0].somModel.sram_dat[2][638][0]=96'h33a608;
sos_loop[0].somModel.sram_ptr[2][638]=2;
sos_loop[0].somModel.sram_dat[2][639][0]=96'h291e21;
sos_loop[0].somModel.sram_ptr[2][639]=2;
sos_loop[0].somModel.sram_dat[2][640][0]=96'hc4dc56;
sos_loop[0].somModel.sram_ptr[2][640]=2;
sos_loop[0].somModel.sram_dat[2][641][0]=96'h1b53a4;
sos_loop[0].somModel.sram_ptr[2][641]=2;
sos_loop[0].somModel.sram_dat[2][642][0]=96'h9d22f;
sos_loop[0].somModel.sram_ptr[2][642]=2;
sos_loop[0].somModel.sram_dat[2][643][0]=96'h5a1b8f;
sos_loop[0].somModel.sram_ptr[2][643]=2;
sos_loop[0].somModel.sram_dat[2][644][0]=96'he01679;
sos_loop[0].somModel.sram_ptr[2][644]=2;
sos_loop[0].somModel.sram_dat[2][645][0]=96'h44e0ed;
sos_loop[0].somModel.sram_ptr[2][645]=2;
sos_loop[0].somModel.sram_dat[2][646][0]=96'hc9bb74;
sos_loop[0].somModel.sram_ptr[2][646]=2;
sos_loop[0].somModel.sram_dat[2][647][0]=96'h5c1683;
sos_loop[0].somModel.sram_ptr[2][647]=2;
sos_loop[0].somModel.sram_dat[2][648][0]=96'h5fbc9d;
sos_loop[0].somModel.sram_ptr[2][648]=2;
sos_loop[0].somModel.sram_dat[2][649][0]=96'hbc2b03;
sos_loop[0].somModel.sram_ptr[2][649]=2;
sos_loop[0].somModel.sram_dat[2][650][0]=96'h44df86;
sos_loop[0].somModel.sram_ptr[2][650]=2;
sos_loop[0].somModel.sram_dat[2][651][0]=96'hdadec5;
sos_loop[0].somModel.sram_ptr[2][651]=2;
sos_loop[0].somModel.sram_dat[2][652][0]=96'h2fa3c2;
sos_loop[0].somModel.sram_ptr[2][652]=2;
sos_loop[0].somModel.sram_dat[2][653][0]=96'h795c0b;
sos_loop[0].somModel.sram_ptr[2][653]=2;
sos_loop[0].somModel.sram_dat[2][654][0]=96'hc6f84e;
sos_loop[0].somModel.sram_ptr[2][654]=2;
sos_loop[0].somModel.sram_dat[2][655][0]=96'hb16934;
sos_loop[0].somModel.sram_ptr[2][655]=2;
sos_loop[0].somModel.sram_dat[2][656][0]=96'h9460ec;
sos_loop[0].somModel.sram_ptr[2][656]=2;
sos_loop[0].somModel.sram_dat[2][657][0]=96'h961e88;
sos_loop[0].somModel.sram_ptr[2][657]=2;
sos_loop[0].somModel.sram_dat[2][658][0]=96'hc93603;
sos_loop[0].somModel.sram_ptr[2][658]=2;
sos_loop[0].somModel.sram_dat[2][659][0]=96'hf71bb0;
sos_loop[0].somModel.sram_ptr[2][659]=2;
sos_loop[0].somModel.sram_dat[2][660][0]=96'hb1611c;
sos_loop[0].somModel.sram_ptr[2][660]=2;
sos_loop[0].somModel.sram_dat[2][661][0]=96'hec7932;
sos_loop[0].somModel.sram_ptr[2][661]=2;
sos_loop[0].somModel.sram_dat[2][662][0]=96'h43bb09;
sos_loop[0].somModel.sram_ptr[2][662]=2;
sos_loop[0].somModel.sram_dat[2][663][0]=96'h40cb8;
sos_loop[0].somModel.sram_ptr[2][663]=2;
sos_loop[0].somModel.sram_dat[2][664][0]=96'h85d475;
sos_loop[0].somModel.sram_ptr[2][664]=2;
sos_loop[0].somModel.sram_dat[2][665][0]=96'ha661a8;
sos_loop[0].somModel.sram_ptr[2][665]=2;
sos_loop[0].somModel.sram_dat[2][666][0]=96'hf38b5;
sos_loop[0].somModel.sram_ptr[2][666]=2;
sos_loop[0].somModel.sram_dat[2][667][0]=96'h986622;
sos_loop[0].somModel.sram_ptr[2][667]=2;
sos_loop[0].somModel.sram_dat[2][668][0]=96'h72876e;
sos_loop[0].somModel.sram_ptr[2][668]=2;
sos_loop[0].somModel.sram_dat[2][669][0]=96'h26c981;
sos_loop[0].somModel.sram_ptr[2][669]=2;
sos_loop[0].somModel.sram_dat[2][670][0]=96'hc3c23a;
sos_loop[0].somModel.sram_ptr[2][670]=2;
sos_loop[0].somModel.sram_dat[2][671][0]=96'h907259;
sos_loop[0].somModel.sram_ptr[2][671]=2;
sos_loop[0].somModel.sram_dat[2][672][0]=96'h52165d;
sos_loop[0].somModel.sram_ptr[2][672]=2;
sos_loop[0].somModel.sram_dat[2][673][0]=96'h95fcd7;
sos_loop[0].somModel.sram_ptr[2][673]=2;
sos_loop[0].somModel.sram_dat[2][674][0]=96'h2dc5de;
sos_loop[0].somModel.sram_ptr[2][674]=2;
sos_loop[0].somModel.sram_dat[2][675][0]=96'h3bd5a3;
sos_loop[0].somModel.sram_ptr[2][675]=2;
sos_loop[0].somModel.sram_dat[2][676][0]=96'ha551ba;
sos_loop[0].somModel.sram_ptr[2][676]=2;
sos_loop[0].somModel.sram_dat[2][677][0]=96'h35e5cb;
sos_loop[0].somModel.sram_ptr[2][677]=2;
sos_loop[0].somModel.sram_dat[2][678][0]=96'hc960bd;
sos_loop[0].somModel.sram_ptr[2][678]=2;
sos_loop[0].somModel.sram_dat[2][679][0]=96'h23b8b6;
sos_loop[0].somModel.sram_ptr[2][679]=2;
sos_loop[0].somModel.sram_dat[2][680][0]=96'hd4d778;
sos_loop[0].somModel.sram_ptr[2][680]=2;
sos_loop[0].somModel.sram_dat[2][681][0]=96'hea3ee3;
sos_loop[0].somModel.sram_ptr[2][681]=2;
sos_loop[0].somModel.sram_dat[2][682][0]=96'h1d84d3;
sos_loop[0].somModel.sram_ptr[2][682]=2;
sos_loop[0].somModel.sram_dat[2][683][0]=96'h77135c;
sos_loop[0].somModel.sram_ptr[2][683]=2;
sos_loop[0].somModel.sram_dat[2][684][0]=96'h61df00;
sos_loop[0].somModel.sram_ptr[2][684]=2;
sos_loop[0].somModel.sram_dat[2][685][0]=96'ha9a5bc;
sos_loop[0].somModel.sram_ptr[2][685]=2;
sos_loop[0].somModel.sram_dat[2][686][0]=96'hba4d19;
sos_loop[0].somModel.sram_ptr[2][686]=2;
sos_loop[0].somModel.sram_dat[2][687][0]=96'hccf409;
sos_loop[0].somModel.sram_ptr[2][687]=2;
sos_loop[0].somModel.sram_dat[2][688][0]=96'h85da8d;
sos_loop[0].somModel.sram_ptr[2][688]=2;
sos_loop[0].somModel.sram_dat[2][689][0]=96'h615d80;
sos_loop[0].somModel.sram_ptr[2][689]=2;
sos_loop[0].somModel.sram_dat[2][690][0]=96'h726469;
sos_loop[0].somModel.sram_ptr[2][690]=2;
sos_loop[0].somModel.sram_dat[2][691][0]=96'h69cc0a;
sos_loop[0].somModel.sram_ptr[2][691]=2;
sos_loop[0].somModel.sram_dat[2][692][0]=96'hb23db7;
sos_loop[0].somModel.sram_ptr[2][692]=2;
sos_loop[0].somModel.sram_dat[2][693][0]=96'h512c45;
sos_loop[0].somModel.sram_ptr[2][693]=2;
sos_loop[0].somModel.sram_dat[2][694][0]=96'hdcffc3;
sos_loop[0].somModel.sram_ptr[2][694]=2;
sos_loop[0].somModel.sram_dat[2][695][0]=96'hcc8fd4;
sos_loop[0].somModel.sram_ptr[2][695]=2;
sos_loop[0].somModel.sram_dat[2][696][0]=96'hac910e;
sos_loop[0].somModel.sram_ptr[2][696]=2;
sos_loop[0].somModel.sram_dat[2][697][0]=96'h66efed;
sos_loop[0].somModel.sram_ptr[2][697]=2;
sos_loop[0].somModel.sram_dat[2][698][0]=96'hd0094e;
sos_loop[0].somModel.sram_ptr[2][698]=2;
sos_loop[0].somModel.sram_dat[2][699][0]=96'hc23370;
sos_loop[0].somModel.sram_ptr[2][699]=2;
sos_loop[0].somModel.sram_dat[2][700][0]=96'hace597;
sos_loop[0].somModel.sram_ptr[2][700]=2;
sos_loop[0].somModel.cfg_tbl_sel[2] = 2;
sos_loop[0].somModel.cfg_dat_sel[2] = 0;
sos_loop[0].somModel.cfg_dat_vld[2] = 1;
sos_loop[0].somModel.cfg_miss_ptr[2] = 0;
sos_loop[0].somModel.tcam_data[3][0][0]=80'h00000000000000000000;
sos_loop[0].somModel.tcam_mask[3][0][0]=80'hffffffffffffffffffff;
sos_loop[0].somModel.tcam_data[3][1][0]=80'h0000000000000093d46a;
sos_loop[0].somModel.tcam_mask[3][1][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][2][0]=80'h00000000000000d2356f;
sos_loop[0].somModel.tcam_mask[3][2][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][3][0]=80'h00000000000000676259;
sos_loop[0].somModel.tcam_mask[3][3][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][4][0]=80'h0000000000000046079b;
sos_loop[0].somModel.tcam_mask[3][4][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][5][0]=80'h000000000000008c8892;
sos_loop[0].somModel.tcam_mask[3][5][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][6][0]=80'h0000000000000017cf44;
sos_loop[0].somModel.tcam_mask[3][6][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][7][0]=80'h00000000000000bc724b;
sos_loop[0].somModel.tcam_mask[3][7][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][8][0]=80'h00000000000000e97981;
sos_loop[0].somModel.tcam_mask[3][8][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][9][0]=80'h0000000000000077a9de;
sos_loop[0].somModel.tcam_mask[3][9][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][10][0]=80'h000000000000002b7a6c;
sos_loop[0].somModel.tcam_mask[3][10][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][11][0]=80'h00000000000000504864;
sos_loop[0].somModel.tcam_mask[3][11][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][12][0]=80'h000000000000008c6bb5;
sos_loop[0].somModel.tcam_mask[3][12][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][13][0]=80'h000000000000007afada;
sos_loop[0].somModel.tcam_mask[3][13][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][14][0]=80'h00000000000000cc3650;
sos_loop[0].somModel.tcam_mask[3][14][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][15][0]=80'h0000000000000000dde1;
sos_loop[0].somModel.tcam_mask[3][15][0]=80'hffffffffffffffff0000;
sos_loop[0].somModel.tcam_data[3][16][0]=80'h0000000000000041bae2;
sos_loop[0].somModel.tcam_mask[3][16][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][17][0]=80'h000000000000004b4f80;
sos_loop[0].somModel.tcam_mask[3][17][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][18][0]=80'h00000000000000ccad23;
sos_loop[0].somModel.tcam_mask[3][18][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][19][0]=80'h00000000000000987d18;
sos_loop[0].somModel.tcam_mask[3][19][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][20][0]=80'h00000000000000354214;
sos_loop[0].somModel.tcam_mask[3][20][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][21][0]=80'h000000000000001b5bf0;
sos_loop[0].somModel.tcam_mask[3][21][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][22][0]=80'h00000000000000cfcfe0;
sos_loop[0].somModel.tcam_mask[3][22][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][23][0]=80'h000000000000005dfdd7;
sos_loop[0].somModel.tcam_mask[3][23][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][24][0]=80'h00000000000000f65193;
sos_loop[0].somModel.tcam_mask[3][24][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][25][0]=80'h00000000000000699932;
sos_loop[0].somModel.tcam_mask[3][25][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][26][0]=80'h000000000000003c1356;
sos_loop[0].somModel.tcam_mask[3][26][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][27][0]=80'h00000000000000da35e5;
sos_loop[0].somModel.tcam_mask[3][27][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][28][0]=80'h00000000000000ab08c2;
sos_loop[0].somModel.tcam_mask[3][28][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][29][0]=80'h0000000000000055162c;
sos_loop[0].somModel.tcam_mask[3][29][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][30][0]=80'h0000000000000048ac99;
sos_loop[0].somModel.tcam_mask[3][30][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][31][0]=80'h00000000000000cf2b64;
sos_loop[0].somModel.tcam_mask[3][31][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][32][0]=80'h00000000000000e09d8f;
sos_loop[0].somModel.tcam_mask[3][32][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][33][0]=80'h000000000000001d11e0;
sos_loop[0].somModel.tcam_mask[3][33][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][34][0]=80'h00000000000000dc6d6f;
sos_loop[0].somModel.tcam_mask[3][34][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][35][0]=80'h0000000000000051d87e;
sos_loop[0].somModel.tcam_mask[3][35][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][36][0]=80'h00000000000000a23c19;
sos_loop[0].somModel.tcam_mask[3][36][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][37][0]=80'h00000000000000a8d569;
sos_loop[0].somModel.tcam_mask[3][37][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][38][0]=80'h000000000000009d9ed7;
sos_loop[0].somModel.tcam_mask[3][38][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][39][0]=80'h0000000000000040e4d5;
sos_loop[0].somModel.tcam_mask[3][39][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][40][0]=80'h000000000000006b550f;
sos_loop[0].somModel.tcam_mask[3][40][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][41][0]=80'h00000000000000b29e2e;
sos_loop[0].somModel.tcam_mask[3][41][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][42][0]=80'h000000000000002e7cf1;
sos_loop[0].somModel.tcam_mask[3][42][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][43][0]=80'h000000000000009200e3;
sos_loop[0].somModel.tcam_mask[3][43][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][44][0]=80'h00000000000000d9b933;
sos_loop[0].somModel.tcam_mask[3][44][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][45][0]=80'h00000000000000ed726f;
sos_loop[0].somModel.tcam_mask[3][45][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][46][0]=80'h000000000000005a968d;
sos_loop[0].somModel.tcam_mask[3][46][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][47][0]=80'h00000000000000aa89df;
sos_loop[0].somModel.tcam_mask[3][47][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][48][0]=80'h00000000000000c1a0ac;
sos_loop[0].somModel.tcam_mask[3][48][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][49][0]=80'h00000000000000281727;
sos_loop[0].somModel.tcam_mask[3][49][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][50][0]=80'h00000000000000fe964b;
sos_loop[0].somModel.tcam_mask[3][50][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][51][0]=80'h00000000000000649d6a;
sos_loop[0].somModel.tcam_mask[3][51][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][52][0]=80'h00000000000000b66d0f;
sos_loop[0].somModel.tcam_mask[3][52][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][53][0]=80'h00000000000000a77176;
sos_loop[0].somModel.tcam_mask[3][53][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][54][0]=80'h00000000000000ab9e57;
sos_loop[0].somModel.tcam_mask[3][54][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][55][0]=80'h00000000000000e15190;
sos_loop[0].somModel.tcam_mask[3][55][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][56][0]=80'h00000000000000935b3f;
sos_loop[0].somModel.tcam_mask[3][56][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][57][0]=80'h0000000000000007d3e7;
sos_loop[0].somModel.tcam_mask[3][57][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][58][0]=80'h00000000000000d866b3;
sos_loop[0].somModel.tcam_mask[3][58][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][59][0]=80'h000000000000004d2d96;
sos_loop[0].somModel.tcam_mask[3][59][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][60][0]=80'h00000000000000932137;
sos_loop[0].somModel.tcam_mask[3][60][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][61][0]=80'h00000000000000d76cda;
sos_loop[0].somModel.tcam_mask[3][61][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][62][0]=80'h00000000000000cfb810;
sos_loop[0].somModel.tcam_mask[3][62][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][63][0]=80'h000000000000001f5e6f;
sos_loop[0].somModel.tcam_mask[3][63][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][64][0]=80'h000000000000000866e5;
sos_loop[0].somModel.tcam_mask[3][64][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][65][0]=80'h00000000000000552409;
sos_loop[0].somModel.tcam_mask[3][65][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][66][0]=80'h0000000000000006819a;
sos_loop[0].somModel.tcam_mask[3][66][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][67][0]=80'h00000000000000dabaa8;
sos_loop[0].somModel.tcam_mask[3][67][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][68][0]=80'h000000000000002fc8a9;
sos_loop[0].somModel.tcam_mask[3][68][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][69][0]=80'h000000000000005014e0;
sos_loop[0].somModel.tcam_mask[3][69][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][70][0]=80'h00000000000000cc782f;
sos_loop[0].somModel.tcam_mask[3][70][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][71][0]=80'h000000000000006dae2a;
sos_loop[0].somModel.tcam_mask[3][71][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][72][0]=80'h0000000000000039b496;
sos_loop[0].somModel.tcam_mask[3][72][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][73][0]=80'h000000000000001cae91;
sos_loop[0].somModel.tcam_mask[3][73][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][74][0]=80'h00000000000000caff50;
sos_loop[0].somModel.tcam_mask[3][74][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][75][0]=80'h00000000000000033bd4;
sos_loop[0].somModel.tcam_mask[3][75][0]=80'hfffffffffffffffc0000;
sos_loop[0].somModel.tcam_data[3][76][0]=80'h000000000000004cb006;
sos_loop[0].somModel.tcam_mask[3][76][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][77][0]=80'h00000000000000a72599;
sos_loop[0].somModel.tcam_mask[3][77][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][78][0]=80'h0000000000000019efb1;
sos_loop[0].somModel.tcam_mask[3][78][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][79][0]=80'h00000000000000bc0688;
sos_loop[0].somModel.tcam_mask[3][79][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][80][0]=80'h0000000000000037cb96;
sos_loop[0].somModel.tcam_mask[3][80][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][81][0]=80'h0000000000000065d77e;
sos_loop[0].somModel.tcam_mask[3][81][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][82][0]=80'h00000000000000a4e182;
sos_loop[0].somModel.tcam_mask[3][82][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][83][0]=80'h00000000000000f9664b;
sos_loop[0].somModel.tcam_mask[3][83][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][84][0]=80'h00000000000000d9d504;
sos_loop[0].somModel.tcam_mask[3][84][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][85][0]=80'h00000000000000ac6429;
sos_loop[0].somModel.tcam_mask[3][85][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][86][0]=80'h000000000000000587b1;
sos_loop[0].somModel.tcam_mask[3][86][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][87][0]=80'h0000000000000070b9ff;
sos_loop[0].somModel.tcam_mask[3][87][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][88][0]=80'h000000000000007817b3;
sos_loop[0].somModel.tcam_mask[3][88][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][89][0]=80'h000000000000005309c8;
sos_loop[0].somModel.tcam_mask[3][89][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][90][0]=80'h00000000000000263667;
sos_loop[0].somModel.tcam_mask[3][90][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][91][0]=80'h00000000000000baef4d;
sos_loop[0].somModel.tcam_mask[3][91][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][92][0]=80'h000000000000009fe398;
sos_loop[0].somModel.tcam_mask[3][92][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][93][0]=80'h00000000000000f404b2;
sos_loop[0].somModel.tcam_mask[3][93][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][94][0]=80'h00000000000000e66811;
sos_loop[0].somModel.tcam_mask[3][94][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][95][0]=80'h000000000000006c4854;
sos_loop[0].somModel.tcam_mask[3][95][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][96][0]=80'h00000000000000e41fbe;
sos_loop[0].somModel.tcam_mask[3][96][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][97][0]=80'h00000000000000ae926c;
sos_loop[0].somModel.tcam_mask[3][97][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][98][0]=80'h000000000000008b4995;
sos_loop[0].somModel.tcam_mask[3][98][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][99][0]=80'h00000000000000ad9ee1;
sos_loop[0].somModel.tcam_mask[3][99][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][100][0]=80'h00000000000000e9cab6;
sos_loop[0].somModel.tcam_mask[3][100][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][101][0]=80'h00000000000000190690;
sos_loop[0].somModel.tcam_mask[3][101][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][102][0]=80'h00000000000000644cd1;
sos_loop[0].somModel.tcam_mask[3][102][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][103][0]=80'h00000000000000193143;
sos_loop[0].somModel.tcam_mask[3][103][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][104][0]=80'h00000000000000b38da9;
sos_loop[0].somModel.tcam_mask[3][104][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][105][0]=80'h00000000000000ad42fb;
sos_loop[0].somModel.tcam_mask[3][105][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][106][0]=80'h00000000000000f0c8e9;
sos_loop[0].somModel.tcam_mask[3][106][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][107][0]=80'h00000000000000c63e22;
sos_loop[0].somModel.tcam_mask[3][107][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][108][0]=80'h00000000000000ceae4f;
sos_loop[0].somModel.tcam_mask[3][108][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][109][0]=80'h0000000000000081fce1;
sos_loop[0].somModel.tcam_mask[3][109][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][110][0]=80'h000000000000006c8b8a;
sos_loop[0].somModel.tcam_mask[3][110][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][111][0]=80'h00000000000000c9c607;
sos_loop[0].somModel.tcam_mask[3][111][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][112][0]=80'h0000000000000084f36d;
sos_loop[0].somModel.tcam_mask[3][112][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][113][0]=80'h00000000000000476c8a;
sos_loop[0].somModel.tcam_mask[3][113][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][114][0]=80'h00000000000000d0a28d;
sos_loop[0].somModel.tcam_mask[3][114][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][115][0]=80'h00000000000000a88374;
sos_loop[0].somModel.tcam_mask[3][115][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][116][0]=80'h00000000000000ec0149;
sos_loop[0].somModel.tcam_mask[3][116][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][117][0]=80'h00000000000000d54c20;
sos_loop[0].somModel.tcam_mask[3][117][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][118][0]=80'h00000000000000990140;
sos_loop[0].somModel.tcam_mask[3][118][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][119][0]=80'h00000000000000d8c32b;
sos_loop[0].somModel.tcam_mask[3][119][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][120][0]=80'h000000000000009db7f1;
sos_loop[0].somModel.tcam_mask[3][120][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][121][0]=80'h000000000000004fa872;
sos_loop[0].somModel.tcam_mask[3][121][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][122][0]=80'h00000000000000fa834c;
sos_loop[0].somModel.tcam_mask[3][122][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][123][0]=80'h00000000000000640129;
sos_loop[0].somModel.tcam_mask[3][123][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][124][0]=80'h00000000000000472ab0;
sos_loop[0].somModel.tcam_mask[3][124][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][125][0]=80'h00000000000000de8fce;
sos_loop[0].somModel.tcam_mask[3][125][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][126][0]=80'h00000000000000e5dd77;
sos_loop[0].somModel.tcam_mask[3][126][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][127][0]=80'h00000000000000e2e528;
sos_loop[0].somModel.tcam_mask[3][127][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][128][0]=80'h00000000000000c4a88f;
sos_loop[0].somModel.tcam_mask[3][128][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][129][0]=80'h0000000000000036d132;
sos_loop[0].somModel.tcam_mask[3][129][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][130][0]=80'h00000000000000103330;
sos_loop[0].somModel.tcam_mask[3][130][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][131][0]=80'h00000000000000210b4b;
sos_loop[0].somModel.tcam_mask[3][131][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][132][0]=80'h0000000000000023a29c;
sos_loop[0].somModel.tcam_mask[3][132][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][133][0]=80'h0000000000000018d134;
sos_loop[0].somModel.tcam_mask[3][133][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][134][0]=80'h00000000000000902d86;
sos_loop[0].somModel.tcam_mask[3][134][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][135][0]=80'h00000000000000599e1e;
sos_loop[0].somModel.tcam_mask[3][135][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][136][0]=80'h000000000000008b80f3;
sos_loop[0].somModel.tcam_mask[3][136][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][137][0]=80'h00000000000000fdd6d9;
sos_loop[0].somModel.tcam_mask[3][137][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][138][0]=80'h00000000000000a822ed;
sos_loop[0].somModel.tcam_mask[3][138][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][139][0]=80'h00000000000000325c6b;
sos_loop[0].somModel.tcam_mask[3][139][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][140][0]=80'h00000000000000f3a0f1;
sos_loop[0].somModel.tcam_mask[3][140][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][141][0]=80'h0000000000000040625f;
sos_loop[0].somModel.tcam_mask[3][141][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][142][0]=80'h00000000000000062576;
sos_loop[0].somModel.tcam_mask[3][142][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][143][0]=80'h00000000000000247741;
sos_loop[0].somModel.tcam_mask[3][143][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][144][0]=80'h00000000000000e66076;
sos_loop[0].somModel.tcam_mask[3][144][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][145][0]=80'h00000000000000a1bfdb;
sos_loop[0].somModel.tcam_mask[3][145][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][146][0]=80'h00000000000000733a59;
sos_loop[0].somModel.tcam_mask[3][146][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][147][0]=80'h00000000000000d5364d;
sos_loop[0].somModel.tcam_mask[3][147][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][148][0]=80'h00000000000000bf32c7;
sos_loop[0].somModel.tcam_mask[3][148][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][149][0]=80'h00000000000000dc5dbf;
sos_loop[0].somModel.tcam_mask[3][149][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][150][0]=80'h000000000000009a93fb;
sos_loop[0].somModel.tcam_mask[3][150][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][151][0]=80'h00000000000000cf1ba8;
sos_loop[0].somModel.tcam_mask[3][151][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][152][0]=80'h000000000000002a29f0;
sos_loop[0].somModel.tcam_mask[3][152][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][153][0]=80'h00000000000000dbde8b;
sos_loop[0].somModel.tcam_mask[3][153][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][154][0]=80'h00000000000000009fe4;
sos_loop[0].somModel.tcam_mask[3][154][0]=80'hffffffffffffffff0000;
sos_loop[0].somModel.tcam_data[3][155][0]=80'h00000000000000180c0a;
sos_loop[0].somModel.tcam_mask[3][155][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][156][0]=80'h0000000000000088f835;
sos_loop[0].somModel.tcam_mask[3][156][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][157][0]=80'h0000000000000017109f;
sos_loop[0].somModel.tcam_mask[3][157][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][158][0]=80'h00000000000000889713;
sos_loop[0].somModel.tcam_mask[3][158][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][159][0]=80'h0000000000000041b6b6;
sos_loop[0].somModel.tcam_mask[3][159][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][160][0]=80'h00000000000000864de9;
sos_loop[0].somModel.tcam_mask[3][160][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][161][0]=80'h0000000000000007abce;
sos_loop[0].somModel.tcam_mask[3][161][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][162][0]=80'h00000000000000e12c35;
sos_loop[0].somModel.tcam_mask[3][162][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][163][0]=80'h00000000000000301447;
sos_loop[0].somModel.tcam_mask[3][163][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][164][0]=80'h00000000000000076b32;
sos_loop[0].somModel.tcam_mask[3][164][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][165][0]=80'h000000000000004b21b3;
sos_loop[0].somModel.tcam_mask[3][165][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][166][0]=80'h00000000000000a87adb;
sos_loop[0].somModel.tcam_mask[3][166][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][167][0]=80'h000000000000008e26bd;
sos_loop[0].somModel.tcam_mask[3][167][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][168][0]=80'h00000000000000e69464;
sos_loop[0].somModel.tcam_mask[3][168][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][169][0]=80'h00000000000000f1ae69;
sos_loop[0].somModel.tcam_mask[3][169][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][170][0]=80'h000000000000003aec7a;
sos_loop[0].somModel.tcam_mask[3][170][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][171][0]=80'h00000000000000ee62e2;
sos_loop[0].somModel.tcam_mask[3][171][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][172][0]=80'h00000000000000e8bc68;
sos_loop[0].somModel.tcam_mask[3][172][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][173][0]=80'h000000000000005b86a9;
sos_loop[0].somModel.tcam_mask[3][173][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][174][0]=80'h000000000000007871a5;
sos_loop[0].somModel.tcam_mask[3][174][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][175][0]=80'h0000000000000055f1d9;
sos_loop[0].somModel.tcam_mask[3][175][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][176][0]=80'h0000000000000096e694;
sos_loop[0].somModel.tcam_mask[3][176][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][177][0]=80'h000000000000001fe63b;
sos_loop[0].somModel.tcam_mask[3][177][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][178][0]=80'h00000000000000806547;
sos_loop[0].somModel.tcam_mask[3][178][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][179][0]=80'h0000000000000025c72f;
sos_loop[0].somModel.tcam_mask[3][179][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][180][0]=80'h00000000000000a62af6;
sos_loop[0].somModel.tcam_mask[3][180][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][181][0]=80'h000000000000009d5417;
sos_loop[0].somModel.tcam_mask[3][181][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][182][0]=80'h000000000000002c51af;
sos_loop[0].somModel.tcam_mask[3][182][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][183][0]=80'h000000000000002f7ca4;
sos_loop[0].somModel.tcam_mask[3][183][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][184][0]=80'h00000000000000c3d2cf;
sos_loop[0].somModel.tcam_mask[3][184][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][185][0]=80'h000000000000002f8d88;
sos_loop[0].somModel.tcam_mask[3][185][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][186][0]=80'h00000000000000128302;
sos_loop[0].somModel.tcam_mask[3][186][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][187][0]=80'h000000000000003cc6e7;
sos_loop[0].somModel.tcam_mask[3][187][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][188][0]=80'h00000000000000bebdfb;
sos_loop[0].somModel.tcam_mask[3][188][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][189][0]=80'h00000000000000aaacbb;
sos_loop[0].somModel.tcam_mask[3][189][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][190][0]=80'h0000000000000035afca;
sos_loop[0].somModel.tcam_mask[3][190][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][191][0]=80'h000000000000003f635d;
sos_loop[0].somModel.tcam_mask[3][191][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][192][0]=80'h000000000000009dc27f;
sos_loop[0].somModel.tcam_mask[3][192][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][193][0]=80'h00000000000000f64438;
sos_loop[0].somModel.tcam_mask[3][193][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][194][0]=80'h000000000000001cde19;
sos_loop[0].somModel.tcam_mask[3][194][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][195][0]=80'h00000000000000ad0b70;
sos_loop[0].somModel.tcam_mask[3][195][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][196][0]=80'h00000000000000b2a22c;
sos_loop[0].somModel.tcam_mask[3][196][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][197][0]=80'h00000000000000c40815;
sos_loop[0].somModel.tcam_mask[3][197][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][198][0]=80'h00000000000000a08a15;
sos_loop[0].somModel.tcam_mask[3][198][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][199][0]=80'h00000000000000294352;
sos_loop[0].somModel.tcam_mask[3][199][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][200][0]=80'h0000000000000009f922;
sos_loop[0].somModel.tcam_mask[3][200][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][201][0]=80'h00000000000000c44933;
sos_loop[0].somModel.tcam_mask[3][201][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][202][0]=80'h00000000000000cba9fb;
sos_loop[0].somModel.tcam_mask[3][202][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][203][0]=80'h00000000000000cee397;
sos_loop[0].somModel.tcam_mask[3][203][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][204][0]=80'h000000000000005ab855;
sos_loop[0].somModel.tcam_mask[3][204][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][205][0]=80'h00000000000000c37cff;
sos_loop[0].somModel.tcam_mask[3][205][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][206][0]=80'h000000000000000f1815;
sos_loop[0].somModel.tcam_mask[3][206][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][207][0]=80'h000000000000001fecf8;
sos_loop[0].somModel.tcam_mask[3][207][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][208][0]=80'h000000000000002f0cd3;
sos_loop[0].somModel.tcam_mask[3][208][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][209][0]=80'h00000000000000cdfdc7;
sos_loop[0].somModel.tcam_mask[3][209][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][210][0]=80'h00000000000000eada3f;
sos_loop[0].somModel.tcam_mask[3][210][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][211][0]=80'h00000000000000c5239f;
sos_loop[0].somModel.tcam_mask[3][211][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][212][0]=80'h000000000000002e0306;
sos_loop[0].somModel.tcam_mask[3][212][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][213][0]=80'h000000000000009b50e8;
sos_loop[0].somModel.tcam_mask[3][213][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][214][0]=80'h00000000000000244d2d;
sos_loop[0].somModel.tcam_mask[3][214][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][215][0]=80'h00000000000000d04cf1;
sos_loop[0].somModel.tcam_mask[3][215][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][216][0]=80'h0000000000000012056a;
sos_loop[0].somModel.tcam_mask[3][216][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][217][0]=80'h0000000000000017ca62;
sos_loop[0].somModel.tcam_mask[3][217][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][218][0]=80'h000000000000003f7a75;
sos_loop[0].somModel.tcam_mask[3][218][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][219][0]=80'h000000000000007a839f;
sos_loop[0].somModel.tcam_mask[3][219][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][220][0]=80'h000000000000000488d5;
sos_loop[0].somModel.tcam_mask[3][220][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][221][0]=80'h0000000000000034ae81;
sos_loop[0].somModel.tcam_mask[3][221][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][222][0]=80'h000000000000001ee202;
sos_loop[0].somModel.tcam_mask[3][222][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][223][0]=80'h00000000000000183ea5;
sos_loop[0].somModel.tcam_mask[3][223][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][224][0]=80'h00000000000000c5cf43;
sos_loop[0].somModel.tcam_mask[3][224][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][225][0]=80'h00000000000000e2bc13;
sos_loop[0].somModel.tcam_mask[3][225][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][226][0]=80'h000000000000001fd051;
sos_loop[0].somModel.tcam_mask[3][226][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][227][0]=80'h000000000000001d970f;
sos_loop[0].somModel.tcam_mask[3][227][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][228][0]=80'h00000000000000c403c7;
sos_loop[0].somModel.tcam_mask[3][228][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][229][0]=80'h0000000000000088f8af;
sos_loop[0].somModel.tcam_mask[3][229][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][230][0]=80'h00000000000000522f39;
sos_loop[0].somModel.tcam_mask[3][230][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][231][0]=80'h00000000000000f385d1;
sos_loop[0].somModel.tcam_mask[3][231][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][232][0]=80'h000000000000009777c8;
sos_loop[0].somModel.tcam_mask[3][232][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][233][0]=80'h00000000000000ffee98;
sos_loop[0].somModel.tcam_mask[3][233][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][234][0]=80'h000000000000008f8852;
sos_loop[0].somModel.tcam_mask[3][234][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][235][0]=80'h0000000000000022a823;
sos_loop[0].somModel.tcam_mask[3][235][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][236][0]=80'h00000000000000aabbdd;
sos_loop[0].somModel.tcam_mask[3][236][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][237][0]=80'h00000000000000c4d792;
sos_loop[0].somModel.tcam_mask[3][237][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][238][0]=80'h000000000000001af82d;
sos_loop[0].somModel.tcam_mask[3][238][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][239][0]=80'h0000000000000012e62a;
sos_loop[0].somModel.tcam_mask[3][239][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][240][0]=80'h0000000000000084feb8;
sos_loop[0].somModel.tcam_mask[3][240][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][241][0]=80'h00000000000000e90935;
sos_loop[0].somModel.tcam_mask[3][241][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][242][0]=80'h00000000000000daeacf;
sos_loop[0].somModel.tcam_mask[3][242][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][243][0]=80'h00000000000000f7fb36;
sos_loop[0].somModel.tcam_mask[3][243][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][244][0]=80'h000000000000000b754c;
sos_loop[0].somModel.tcam_mask[3][244][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][245][0]=80'h0000000000000072a0d2;
sos_loop[0].somModel.tcam_mask[3][245][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][246][0]=80'h0000000000000014c7a8;
sos_loop[0].somModel.tcam_mask[3][246][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][247][0]=80'h000000000000002e7ccb;
sos_loop[0].somModel.tcam_mask[3][247][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][248][0]=80'h00000000000000172d6b;
sos_loop[0].somModel.tcam_mask[3][248][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][249][0]=80'h000000000000005cbd69;
sos_loop[0].somModel.tcam_mask[3][249][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][250][0]=80'h00000000000000838848;
sos_loop[0].somModel.tcam_mask[3][250][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][251][0]=80'h00000000000000e57f48;
sos_loop[0].somModel.tcam_mask[3][251][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][252][0]=80'h00000000000000879954;
sos_loop[0].somModel.tcam_mask[3][252][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][253][0]=80'h000000000000003f3b48;
sos_loop[0].somModel.tcam_mask[3][253][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][254][0]=80'h00000000000000aa15a1;
sos_loop[0].somModel.tcam_mask[3][254][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][255][0]=80'h0000000000000072e889;
sos_loop[0].somModel.tcam_mask[3][255][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][256][0]=80'h0000000000000001b542;
sos_loop[0].somModel.tcam_mask[3][256][0]=80'hfffffffffffffffe0000;
sos_loop[0].somModel.tcam_data[3][257][0]=80'h00000000000000296632;
sos_loop[0].somModel.tcam_mask[3][257][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][258][0]=80'h0000000000000038ad9e;
sos_loop[0].somModel.tcam_mask[3][258][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][259][0]=80'h00000000000000dd5b20;
sos_loop[0].somModel.tcam_mask[3][259][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][260][0]=80'h000000000000007e3d3f;
sos_loop[0].somModel.tcam_mask[3][260][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][261][0]=80'h00000000000000de577e;
sos_loop[0].somModel.tcam_mask[3][261][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][262][0]=80'h000000000000005f90c0;
sos_loop[0].somModel.tcam_mask[3][262][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][263][0]=80'h00000000000000d30cb2;
sos_loop[0].somModel.tcam_mask[3][263][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][264][0]=80'h000000000000008ebe76;
sos_loop[0].somModel.tcam_mask[3][264][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][265][0]=80'h000000000000002d1e33;
sos_loop[0].somModel.tcam_mask[3][265][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][266][0]=80'h0000000000000078e2fd;
sos_loop[0].somModel.tcam_mask[3][266][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][267][0]=80'h000000000000008595a0;
sos_loop[0].somModel.tcam_mask[3][267][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][268][0]=80'h000000000000004d7b60;
sos_loop[0].somModel.tcam_mask[3][268][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][269][0]=80'h000000000000000a5d4d;
sos_loop[0].somModel.tcam_mask[3][269][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][270][0]=80'h00000000000000b6a7b0;
sos_loop[0].somModel.tcam_mask[3][270][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][271][0]=80'h00000000000000b9d0d8;
sos_loop[0].somModel.tcam_mask[3][271][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][272][0]=80'h000000000000007c54d0;
sos_loop[0].somModel.tcam_mask[3][272][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][273][0]=80'h00000000000000000fab;
sos_loop[0].somModel.tcam_mask[3][273][0]=80'hfffffffffffffffff000;
sos_loop[0].somModel.tcam_data[3][274][0]=80'h00000000000000526452;
sos_loop[0].somModel.tcam_mask[3][274][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][275][0]=80'h00000000000000eea715;
sos_loop[0].somModel.tcam_mask[3][275][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][276][0]=80'h00000000000000b958bc;
sos_loop[0].somModel.tcam_mask[3][276][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][277][0]=80'h00000000000000a9b50c;
sos_loop[0].somModel.tcam_mask[3][277][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][278][0]=80'h00000000000000fcbf5c;
sos_loop[0].somModel.tcam_mask[3][278][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][279][0]=80'h00000000000000d7128e;
sos_loop[0].somModel.tcam_mask[3][279][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][280][0]=80'h00000000000000287b14;
sos_loop[0].somModel.tcam_mask[3][280][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][281][0]=80'h0000000000000099d893;
sos_loop[0].somModel.tcam_mask[3][281][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][282][0]=80'h00000000000000ce1be7;
sos_loop[0].somModel.tcam_mask[3][282][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][283][0]=80'h00000000000000275c14;
sos_loop[0].somModel.tcam_mask[3][283][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][284][0]=80'h00000000000000b2ecf6;
sos_loop[0].somModel.tcam_mask[3][284][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][285][0]=80'h0000000000000032209f;
sos_loop[0].somModel.tcam_mask[3][285][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][286][0]=80'h000000000000008890e9;
sos_loop[0].somModel.tcam_mask[3][286][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][287][0]=80'h000000000000005df3a2;
sos_loop[0].somModel.tcam_mask[3][287][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][288][0]=80'h00000000000000681f7e;
sos_loop[0].somModel.tcam_mask[3][288][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][289][0]=80'h0000000000000052ac42;
sos_loop[0].somModel.tcam_mask[3][289][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][290][0]=80'h0000000000000062b76d;
sos_loop[0].somModel.tcam_mask[3][290][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][291][0]=80'h000000000000002a3054;
sos_loop[0].somModel.tcam_mask[3][291][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][292][0]=80'h00000000000000a6aacb;
sos_loop[0].somModel.tcam_mask[3][292][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][293][0]=80'h00000000000000fad7b0;
sos_loop[0].somModel.tcam_mask[3][293][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][294][0]=80'h00000000000000e45af7;
sos_loop[0].somModel.tcam_mask[3][294][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][295][0]=80'h000000000000001b8312;
sos_loop[0].somModel.tcam_mask[3][295][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][296][0]=80'h000000000000004d7686;
sos_loop[0].somModel.tcam_mask[3][296][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][297][0]=80'h000000000000009e9f11;
sos_loop[0].somModel.tcam_mask[3][297][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][298][0]=80'h000000000000003752b8;
sos_loop[0].somModel.tcam_mask[3][298][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][299][0]=80'h000000000000009fff19;
sos_loop[0].somModel.tcam_mask[3][299][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][300][0]=80'h000000000000003deeb0;
sos_loop[0].somModel.tcam_mask[3][300][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][301][0]=80'h000000000000004d0cc0;
sos_loop[0].somModel.tcam_mask[3][301][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][302][0]=80'h00000000000000ad4e0b;
sos_loop[0].somModel.tcam_mask[3][302][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][303][0]=80'h00000000000000d93c76;
sos_loop[0].somModel.tcam_mask[3][303][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][304][0]=80'h00000000000000a363f3;
sos_loop[0].somModel.tcam_mask[3][304][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][305][0]=80'h00000000000000fe7a4a;
sos_loop[0].somModel.tcam_mask[3][305][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][306][0]=80'h000000000000006750fd;
sos_loop[0].somModel.tcam_mask[3][306][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][307][0]=80'h00000000000000fa4199;
sos_loop[0].somModel.tcam_mask[3][307][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][308][0]=80'h00000000000000d91f85;
sos_loop[0].somModel.tcam_mask[3][308][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][309][0]=80'h000000000000006021c5;
sos_loop[0].somModel.tcam_mask[3][309][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][310][0]=80'h00000000000000b7fc65;
sos_loop[0].somModel.tcam_mask[3][310][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][311][0]=80'h000000000000000d6e41;
sos_loop[0].somModel.tcam_mask[3][311][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][312][0]=80'h000000000000001fc6a1;
sos_loop[0].somModel.tcam_mask[3][312][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][313][0]=80'h00000000000000d152b0;
sos_loop[0].somModel.tcam_mask[3][313][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][314][0]=80'h000000000000002f8780;
sos_loop[0].somModel.tcam_mask[3][314][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][315][0]=80'h000000000000000a9948;
sos_loop[0].somModel.tcam_mask[3][315][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][316][0]=80'h00000000000000249ab8;
sos_loop[0].somModel.tcam_mask[3][316][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][317][0]=80'h00000000000000472875;
sos_loop[0].somModel.tcam_mask[3][317][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][318][0]=80'h000000000000006d2196;
sos_loop[0].somModel.tcam_mask[3][318][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][319][0]=80'h0000000000000010373f;
sos_loop[0].somModel.tcam_mask[3][319][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][320][0]=80'h00000000000000c0f50e;
sos_loop[0].somModel.tcam_mask[3][320][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][321][0]=80'h00000000000000dd84a8;
sos_loop[0].somModel.tcam_mask[3][321][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][322][0]=80'h00000000000000324444;
sos_loop[0].somModel.tcam_mask[3][322][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][323][0]=80'h00000000000000b11fe3;
sos_loop[0].somModel.tcam_mask[3][323][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][324][0]=80'h00000000000000d3c003;
sos_loop[0].somModel.tcam_mask[3][324][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][325][0]=80'h0000000000000022c068;
sos_loop[0].somModel.tcam_mask[3][325][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][326][0]=80'h00000000000000200557;
sos_loop[0].somModel.tcam_mask[3][326][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][327][0]=80'h00000000000000d760d5;
sos_loop[0].somModel.tcam_mask[3][327][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][328][0]=80'h00000000000000404d84;
sos_loop[0].somModel.tcam_mask[3][328][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][329][0]=80'h0000000000000038a6a0;
sos_loop[0].somModel.tcam_mask[3][329][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][330][0]=80'h000000000000003a4640;
sos_loop[0].somModel.tcam_mask[3][330][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][331][0]=80'h000000000000004a10b1;
sos_loop[0].somModel.tcam_mask[3][331][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][332][0]=80'h00000000000000b30115;
sos_loop[0].somModel.tcam_mask[3][332][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][333][0]=80'h000000000000008aeaa5;
sos_loop[0].somModel.tcam_mask[3][333][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][334][0]=80'h00000000000000f1cc59;
sos_loop[0].somModel.tcam_mask[3][334][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][335][0]=80'h000000000000007f6f35;
sos_loop[0].somModel.tcam_mask[3][335][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][336][0]=80'h00000000000000465838;
sos_loop[0].somModel.tcam_mask[3][336][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][337][0]=80'h00000000000000c08db5;
sos_loop[0].somModel.tcam_mask[3][337][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][338][0]=80'h00000000000000fd7be1;
sos_loop[0].somModel.tcam_mask[3][338][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][339][0]=80'h0000000000000000a0f3;
sos_loop[0].somModel.tcam_mask[3][339][0]=80'hffffffffffffffff0000;
sos_loop[0].somModel.tcam_data[3][340][0]=80'h00000000000000b91869;
sos_loop[0].somModel.tcam_mask[3][340][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][341][0]=80'h00000000000000c0ad63;
sos_loop[0].somModel.tcam_mask[3][341][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][342][0]=80'h00000000000000b08e22;
sos_loop[0].somModel.tcam_mask[3][342][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][343][0]=80'h00000000000000f68553;
sos_loop[0].somModel.tcam_mask[3][343][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][344][0]=80'h0000000000000064927f;
sos_loop[0].somModel.tcam_mask[3][344][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][345][0]=80'h0000000000000083a02e;
sos_loop[0].somModel.tcam_mask[3][345][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][346][0]=80'h00000000000000be5a96;
sos_loop[0].somModel.tcam_mask[3][346][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][347][0]=80'h000000000000006e40d1;
sos_loop[0].somModel.tcam_mask[3][347][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][348][0]=80'h00000000000000f76daa;
sos_loop[0].somModel.tcam_mask[3][348][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][349][0]=80'h00000000000000260806;
sos_loop[0].somModel.tcam_mask[3][349][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][350][0]=80'h00000000000000aaf348;
sos_loop[0].somModel.tcam_mask[3][350][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][351][0]=80'h000000000000000be1a7;
sos_loop[0].somModel.tcam_mask[3][351][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][352][0]=80'h00000000000000a59283;
sos_loop[0].somModel.tcam_mask[3][352][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][353][0]=80'h000000000000009fd1ab;
sos_loop[0].somModel.tcam_mask[3][353][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][354][0]=80'h000000000000008acbff;
sos_loop[0].somModel.tcam_mask[3][354][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][355][0]=80'h000000000000004deca7;
sos_loop[0].somModel.tcam_mask[3][355][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][356][0]=80'h0000000000000028e13a;
sos_loop[0].somModel.tcam_mask[3][356][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][357][0]=80'h00000000000000a299ca;
sos_loop[0].somModel.tcam_mask[3][357][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][358][0]=80'h0000000000000099a477;
sos_loop[0].somModel.tcam_mask[3][358][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][359][0]=80'h0000000000000044a766;
sos_loop[0].somModel.tcam_mask[3][359][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][360][0]=80'h00000000000000d3a394;
sos_loop[0].somModel.tcam_mask[3][360][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][361][0]=80'h00000000000000ecc3e8;
sos_loop[0].somModel.tcam_mask[3][361][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][362][0]=80'h00000000000000ebab0e;
sos_loop[0].somModel.tcam_mask[3][362][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][363][0]=80'h000000000000007f07a0;
sos_loop[0].somModel.tcam_mask[3][363][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][364][0]=80'h000000000000001940da;
sos_loop[0].somModel.tcam_mask[3][364][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][365][0]=80'h00000000000000dd77fd;
sos_loop[0].somModel.tcam_mask[3][365][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][366][0]=80'h0000000000000027a422;
sos_loop[0].somModel.tcam_mask[3][366][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][367][0]=80'h00000000000000e19559;
sos_loop[0].somModel.tcam_mask[3][367][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][368][0]=80'h00000000000000008d63;
sos_loop[0].somModel.tcam_mask[3][368][0]=80'hffffffffffffffff0000;
sos_loop[0].somModel.tcam_data[3][369][0]=80'h0000000000000001193c;
sos_loop[0].somModel.tcam_mask[3][369][0]=80'hfffffffffffffffe0000;
sos_loop[0].somModel.tcam_data[3][370][0]=80'h0000000000000046a7c0;
sos_loop[0].somModel.tcam_mask[3][370][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][371][0]=80'h00000000000000c71745;
sos_loop[0].somModel.tcam_mask[3][371][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][372][0]=80'h00000000000000ee0321;
sos_loop[0].somModel.tcam_mask[3][372][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][373][0]=80'h0000000000000021c943;
sos_loop[0].somModel.tcam_mask[3][373][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][374][0]=80'h000000000000005334c6;
sos_loop[0].somModel.tcam_mask[3][374][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][375][0]=80'h00000000000000cbd414;
sos_loop[0].somModel.tcam_mask[3][375][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][376][0]=80'h00000000000000ab0538;
sos_loop[0].somModel.tcam_mask[3][376][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][377][0]=80'h00000000000000f176c0;
sos_loop[0].somModel.tcam_mask[3][377][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][378][0]=80'h000000000000008512ed;
sos_loop[0].somModel.tcam_mask[3][378][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][379][0]=80'h00000000000000a0128d;
sos_loop[0].somModel.tcam_mask[3][379][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][380][0]=80'h00000000000000db3124;
sos_loop[0].somModel.tcam_mask[3][380][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][381][0]=80'h000000000000003d7888;
sos_loop[0].somModel.tcam_mask[3][381][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][382][0]=80'h0000000000000006f91b;
sos_loop[0].somModel.tcam_mask[3][382][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][383][0]=80'h00000000000000b21e43;
sos_loop[0].somModel.tcam_mask[3][383][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][384][0]=80'h000000000000008de00c;
sos_loop[0].somModel.tcam_mask[3][384][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][385][0]=80'h00000000000000ad6a91;
sos_loop[0].somModel.tcam_mask[3][385][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][386][0]=80'h000000000000009982b5;
sos_loop[0].somModel.tcam_mask[3][386][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][387][0]=80'h00000000000000f936b6;
sos_loop[0].somModel.tcam_mask[3][387][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][388][0]=80'h00000000000000fb8434;
sos_loop[0].somModel.tcam_mask[3][388][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][389][0]=80'h0000000000000061ac31;
sos_loop[0].somModel.tcam_mask[3][389][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][390][0]=80'h00000000000000000d66;
sos_loop[0].somModel.tcam_mask[3][390][0]=80'hfffffffffffffffff000;
sos_loop[0].somModel.tcam_data[3][391][0]=80'h00000000000000cb4d6b;
sos_loop[0].somModel.tcam_mask[3][391][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][392][0]=80'h00000000000000952555;
sos_loop[0].somModel.tcam_mask[3][392][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][393][0]=80'h00000000000000d662de;
sos_loop[0].somModel.tcam_mask[3][393][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][394][0]=80'h00000000000000aa0ea6;
sos_loop[0].somModel.tcam_mask[3][394][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][395][0]=80'h00000000000000ba2e0f;
sos_loop[0].somModel.tcam_mask[3][395][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][396][0]=80'h00000000000000f7491c;
sos_loop[0].somModel.tcam_mask[3][396][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][397][0]=80'h000000000000008d68ee;
sos_loop[0].somModel.tcam_mask[3][397][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][398][0]=80'h00000000000000a366a5;
sos_loop[0].somModel.tcam_mask[3][398][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][399][0]=80'h000000000000007672fe;
sos_loop[0].somModel.tcam_mask[3][399][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][400][0]=80'h000000000000004e0e5b;
sos_loop[0].somModel.tcam_mask[3][400][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][401][0]=80'h00000000000000f69f93;
sos_loop[0].somModel.tcam_mask[3][401][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][402][0]=80'h00000000000000dc64a3;
sos_loop[0].somModel.tcam_mask[3][402][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][403][0]=80'h000000000000003e36d7;
sos_loop[0].somModel.tcam_mask[3][403][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][404][0]=80'h0000000000000020cd14;
sos_loop[0].somModel.tcam_mask[3][404][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][405][0]=80'h00000000000000fd80ee;
sos_loop[0].somModel.tcam_mask[3][405][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][406][0]=80'h0000000000000014a853;
sos_loop[0].somModel.tcam_mask[3][406][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][407][0]=80'h00000000000000d34e71;
sos_loop[0].somModel.tcam_mask[3][407][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][408][0]=80'h000000000000004da43e;
sos_loop[0].somModel.tcam_mask[3][408][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][409][0]=80'h000000000000002dcdd0;
sos_loop[0].somModel.tcam_mask[3][409][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][410][0]=80'h00000000000000ff51e4;
sos_loop[0].somModel.tcam_mask[3][410][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][411][0]=80'h000000000000005e4c3b;
sos_loop[0].somModel.tcam_mask[3][411][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][412][0]=80'h00000000000000919a50;
sos_loop[0].somModel.tcam_mask[3][412][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][413][0]=80'h0000000000000005c6f6;
sos_loop[0].somModel.tcam_mask[3][413][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][414][0]=80'h000000000000004880e1;
sos_loop[0].somModel.tcam_mask[3][414][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][415][0]=80'h00000000000000b52f6e;
sos_loop[0].somModel.tcam_mask[3][415][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][416][0]=80'h000000000000006330f5;
sos_loop[0].somModel.tcam_mask[3][416][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][417][0]=80'h0000000000000087589c;
sos_loop[0].somModel.tcam_mask[3][417][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][418][0]=80'h00000000000000ae87c5;
sos_loop[0].somModel.tcam_mask[3][418][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][419][0]=80'h0000000000000088b591;
sos_loop[0].somModel.tcam_mask[3][419][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][420][0]=80'h00000000000000a9681c;
sos_loop[0].somModel.tcam_mask[3][420][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][421][0]=80'h000000000000005bfe8c;
sos_loop[0].somModel.tcam_mask[3][421][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][422][0]=80'h00000000000000feeabb;
sos_loop[0].somModel.tcam_mask[3][422][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][423][0]=80'h000000000000005bfef3;
sos_loop[0].somModel.tcam_mask[3][423][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][424][0]=80'h00000000000000c439f5;
sos_loop[0].somModel.tcam_mask[3][424][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][425][0]=80'h00000000000000cbb611;
sos_loop[0].somModel.tcam_mask[3][425][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][426][0]=80'h000000000000006bf841;
sos_loop[0].somModel.tcam_mask[3][426][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][427][0]=80'h0000000000000014eb96;
sos_loop[0].somModel.tcam_mask[3][427][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][428][0]=80'h00000000000000cb6ce3;
sos_loop[0].somModel.tcam_mask[3][428][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][429][0]=80'h00000000000000be0907;
sos_loop[0].somModel.tcam_mask[3][429][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][430][0]=80'h00000000000000f515b5;
sos_loop[0].somModel.tcam_mask[3][430][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][431][0]=80'h00000000000000d4b21b;
sos_loop[0].somModel.tcam_mask[3][431][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][432][0]=80'h00000000000000aed1b5;
sos_loop[0].somModel.tcam_mask[3][432][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][433][0]=80'h000000000000000187e1;
sos_loop[0].somModel.tcam_mask[3][433][0]=80'hfffffffffffffffe0000;
sos_loop[0].somModel.tcam_data[3][434][0]=80'h000000000000003bf896;
sos_loop[0].somModel.tcam_mask[3][434][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][435][0]=80'h00000000000000d53055;
sos_loop[0].somModel.tcam_mask[3][435][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][436][0]=80'h00000000000000d85a46;
sos_loop[0].somModel.tcam_mask[3][436][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][437][0]=80'h00000000000000b70da5;
sos_loop[0].somModel.tcam_mask[3][437][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][438][0]=80'h00000000000000f14efb;
sos_loop[0].somModel.tcam_mask[3][438][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][439][0]=80'h00000000000000ceed54;
sos_loop[0].somModel.tcam_mask[3][439][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][440][0]=80'h000000000000001c63cc;
sos_loop[0].somModel.tcam_mask[3][440][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][441][0]=80'h000000000000002e657b;
sos_loop[0].somModel.tcam_mask[3][441][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][442][0]=80'h000000000000001b7bb1;
sos_loop[0].somModel.tcam_mask[3][442][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][443][0]=80'h00000000000000a490bb;
sos_loop[0].somModel.tcam_mask[3][443][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][444][0]=80'h0000000000000077f7c3;
sos_loop[0].somModel.tcam_mask[3][444][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][445][0]=80'h00000000000000ce3879;
sos_loop[0].somModel.tcam_mask[3][445][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][446][0]=80'h000000000000003d62f7;
sos_loop[0].somModel.tcam_mask[3][446][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][447][0]=80'h00000000000000d3c317;
sos_loop[0].somModel.tcam_mask[3][447][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][448][0]=80'h00000000000000cd4052;
sos_loop[0].somModel.tcam_mask[3][448][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][449][0]=80'h00000000000000366029;
sos_loop[0].somModel.tcam_mask[3][449][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][450][0]=80'h00000000000000249c31;
sos_loop[0].somModel.tcam_mask[3][450][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][451][0]=80'h00000000000000f85353;
sos_loop[0].somModel.tcam_mask[3][451][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][452][0]=80'h00000000000000ba861d;
sos_loop[0].somModel.tcam_mask[3][452][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][453][0]=80'h000000000000007b4f14;
sos_loop[0].somModel.tcam_mask[3][453][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][454][0]=80'h00000000000000e9a8b0;
sos_loop[0].somModel.tcam_mask[3][454][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][455][0]=80'h0000000000000048daff;
sos_loop[0].somModel.tcam_mask[3][455][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][456][0]=80'h0000000000000009eeb3;
sos_loop[0].somModel.tcam_mask[3][456][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][457][0]=80'h0000000000000001ea67;
sos_loop[0].somModel.tcam_mask[3][457][0]=80'hfffffffffffffffe0000;
sos_loop[0].somModel.tcam_data[3][458][0]=80'h00000000000000b2c532;
sos_loop[0].somModel.tcam_mask[3][458][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][459][0]=80'h000000000000008cdabd;
sos_loop[0].somModel.tcam_mask[3][459][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][460][0]=80'h00000000000000e33611;
sos_loop[0].somModel.tcam_mask[3][460][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][461][0]=80'h00000000000000888646;
sos_loop[0].somModel.tcam_mask[3][461][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][462][0]=80'h000000000000007532ec;
sos_loop[0].somModel.tcam_mask[3][462][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][463][0]=80'h00000000000000ef77eb;
sos_loop[0].somModel.tcam_mask[3][463][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][464][0]=80'h00000000000000836a74;
sos_loop[0].somModel.tcam_mask[3][464][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][465][0]=80'h0000000000000060abde;
sos_loop[0].somModel.tcam_mask[3][465][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][466][0]=80'h000000000000001fb207;
sos_loop[0].somModel.tcam_mask[3][466][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][467][0]=80'h000000000000001fd4bb;
sos_loop[0].somModel.tcam_mask[3][467][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][468][0]=80'h00000000000000e37673;
sos_loop[0].somModel.tcam_mask[3][468][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][469][0]=80'h00000000000000e78f3e;
sos_loop[0].somModel.tcam_mask[3][469][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][470][0]=80'h00000000000000f089bc;
sos_loop[0].somModel.tcam_mask[3][470][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][471][0]=80'h00000000000000989a46;
sos_loop[0].somModel.tcam_mask[3][471][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][472][0]=80'h0000000000000004872d;
sos_loop[0].somModel.tcam_mask[3][472][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][473][0]=80'h000000000000007d4a59;
sos_loop[0].somModel.tcam_mask[3][473][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][474][0]=80'h0000000000000079148c;
sos_loop[0].somModel.tcam_mask[3][474][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][475][0]=80'h00000000000000ca4d53;
sos_loop[0].somModel.tcam_mask[3][475][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][476][0]=80'h00000000000000318859;
sos_loop[0].somModel.tcam_mask[3][476][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][477][0]=80'h00000000000000d19af7;
sos_loop[0].somModel.tcam_mask[3][477][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][478][0]=80'h00000000000000270545;
sos_loop[0].somModel.tcam_mask[3][478][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][479][0]=80'h0000000000000094a8f5;
sos_loop[0].somModel.tcam_mask[3][479][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][480][0]=80'h00000000000000fd4a65;
sos_loop[0].somModel.tcam_mask[3][480][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][481][0]=80'h0000000000000014a4ed;
sos_loop[0].somModel.tcam_mask[3][481][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][482][0]=80'h00000000000000b279ba;
sos_loop[0].somModel.tcam_mask[3][482][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][483][0]=80'h0000000000000063905b;
sos_loop[0].somModel.tcam_mask[3][483][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][484][0]=80'h00000000000000528285;
sos_loop[0].somModel.tcam_mask[3][484][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][485][0]=80'h00000000000000bd6eb1;
sos_loop[0].somModel.tcam_mask[3][485][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][486][0]=80'h00000000000000136e6c;
sos_loop[0].somModel.tcam_mask[3][486][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][487][0]=80'h000000000000009b3456;
sos_loop[0].somModel.tcam_mask[3][487][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][488][0]=80'h00000000000000254c0a;
sos_loop[0].somModel.tcam_mask[3][488][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][489][0]=80'h00000000000000ec438c;
sos_loop[0].somModel.tcam_mask[3][489][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][490][0]=80'h0000000000000084699d;
sos_loop[0].somModel.tcam_mask[3][490][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][491][0]=80'h000000000000000d0224;
sos_loop[0].somModel.tcam_mask[3][491][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][492][0]=80'h00000000000000c49916;
sos_loop[0].somModel.tcam_mask[3][492][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][493][0]=80'h00000000000000ff4173;
sos_loop[0].somModel.tcam_mask[3][493][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][494][0]=80'h0000000000000081bccf;
sos_loop[0].somModel.tcam_mask[3][494][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][495][0]=80'h000000000000006fed17;
sos_loop[0].somModel.tcam_mask[3][495][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][496][0]=80'h000000000000002329d9;
sos_loop[0].somModel.tcam_mask[3][496][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][497][0]=80'h00000000000000e35295;
sos_loop[0].somModel.tcam_mask[3][497][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][498][0]=80'h0000000000000097a6ce;
sos_loop[0].somModel.tcam_mask[3][498][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][499][0]=80'h000000000000007355fd;
sos_loop[0].somModel.tcam_mask[3][499][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][500][0]=80'h00000000000000b5e794;
sos_loop[0].somModel.tcam_mask[3][500][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][501][0]=80'h000000000000003295ab;
sos_loop[0].somModel.tcam_mask[3][501][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][502][0]=80'h00000000000000eca5ce;
sos_loop[0].somModel.tcam_mask[3][502][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][503][0]=80'h0000000000000087bf14;
sos_loop[0].somModel.tcam_mask[3][503][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][504][0]=80'h00000000000000a166f5;
sos_loop[0].somModel.tcam_mask[3][504][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][505][0]=80'h00000000000000c0b98a;
sos_loop[0].somModel.tcam_mask[3][505][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][506][0]=80'h00000000000000452cdc;
sos_loop[0].somModel.tcam_mask[3][506][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][507][0]=80'h0000000000000078e1e0;
sos_loop[0].somModel.tcam_mask[3][507][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][508][0]=80'h0000000000000092eb8c;
sos_loop[0].somModel.tcam_mask[3][508][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][509][0]=80'h00000000000000129629;
sos_loop[0].somModel.tcam_mask[3][509][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][510][0]=80'h00000000000000bc837b;
sos_loop[0].somModel.tcam_mask[3][510][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][511][0]=80'h000000000000009cda8f;
sos_loop[0].somModel.tcam_mask[3][511][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][512][0]=80'h000000000000003e36f7;
sos_loop[0].somModel.tcam_mask[3][512][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][513][0]=80'h000000000000008a27cd;
sos_loop[0].somModel.tcam_mask[3][513][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][514][0]=80'h00000000000000462c62;
sos_loop[0].somModel.tcam_mask[3][514][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][515][0]=80'h00000000000000dfcade;
sos_loop[0].somModel.tcam_mask[3][515][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][516][0]=80'h000000000000008989c8;
sos_loop[0].somModel.tcam_mask[3][516][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][517][0]=80'h000000000000006c0294;
sos_loop[0].somModel.tcam_mask[3][517][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][518][0]=80'h00000000000000bcd2eb;
sos_loop[0].somModel.tcam_mask[3][518][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][519][0]=80'h000000000000003bff68;
sos_loop[0].somModel.tcam_mask[3][519][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][520][0]=80'h000000000000006b9b27;
sos_loop[0].somModel.tcam_mask[3][520][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][521][0]=80'h0000000000000022b3ea;
sos_loop[0].somModel.tcam_mask[3][521][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][522][0]=80'h0000000000000041688a;
sos_loop[0].somModel.tcam_mask[3][522][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][523][0]=80'h00000000000000e21345;
sos_loop[0].somModel.tcam_mask[3][523][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][524][0]=80'h0000000000000073d32b;
sos_loop[0].somModel.tcam_mask[3][524][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][525][0]=80'h00000000000000a2a953;
sos_loop[0].somModel.tcam_mask[3][525][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][526][0]=80'h000000000000004e430c;
sos_loop[0].somModel.tcam_mask[3][526][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][527][0]=80'h0000000000000064d84c;
sos_loop[0].somModel.tcam_mask[3][527][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][528][0]=80'h000000000000002f0b4c;
sos_loop[0].somModel.tcam_mask[3][528][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][529][0]=80'h000000000000003b69f1;
sos_loop[0].somModel.tcam_mask[3][529][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][530][0]=80'h000000000000000ac0c0;
sos_loop[0].somModel.tcam_mask[3][530][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][531][0]=80'h0000000000000002cb8c;
sos_loop[0].somModel.tcam_mask[3][531][0]=80'hfffffffffffffffc0000;
sos_loop[0].somModel.tcam_data[3][532][0]=80'h00000000000000c8973d;
sos_loop[0].somModel.tcam_mask[3][532][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][533][0]=80'h0000000000000063403b;
sos_loop[0].somModel.tcam_mask[3][533][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][534][0]=80'h000000000000003b10ba;
sos_loop[0].somModel.tcam_mask[3][534][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][535][0]=80'h000000000000002ce7ba;
sos_loop[0].somModel.tcam_mask[3][535][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][536][0]=80'h0000000000000000ea87;
sos_loop[0].somModel.tcam_mask[3][536][0]=80'hffffffffffffffff0000;
sos_loop[0].somModel.tcam_data[3][537][0]=80'h0000000000000050badf;
sos_loop[0].somModel.tcam_mask[3][537][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][538][0]=80'h000000000000005b2fbb;
sos_loop[0].somModel.tcam_mask[3][538][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][539][0]=80'h00000000000000ac32d9;
sos_loop[0].somModel.tcam_mask[3][539][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][540][0]=80'h00000000000000175207;
sos_loop[0].somModel.tcam_mask[3][540][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][541][0]=80'h00000000000000ce27f9;
sos_loop[0].somModel.tcam_mask[3][541][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][542][0]=80'h0000000000000075d740;
sos_loop[0].somModel.tcam_mask[3][542][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][543][0]=80'h0000000000000076d79a;
sos_loop[0].somModel.tcam_mask[3][543][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][544][0]=80'h000000000000007390f8;
sos_loop[0].somModel.tcam_mask[3][544][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][545][0]=80'h00000000000000b963bf;
sos_loop[0].somModel.tcam_mask[3][545][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][546][0]=80'h00000000000000026405;
sos_loop[0].somModel.tcam_mask[3][546][0]=80'hfffffffffffffffc0000;
sos_loop[0].somModel.tcam_data[3][547][0]=80'h00000000000000a04b21;
sos_loop[0].somModel.tcam_mask[3][547][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][548][0]=80'h00000000000000a30541;
sos_loop[0].somModel.tcam_mask[3][548][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][549][0]=80'h000000000000008927b6;
sos_loop[0].somModel.tcam_mask[3][549][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][550][0]=80'h000000000000009cc1c0;
sos_loop[0].somModel.tcam_mask[3][550][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][551][0]=80'h000000000000003ba3f5;
sos_loop[0].somModel.tcam_mask[3][551][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][552][0]=80'h00000000000000352e1d;
sos_loop[0].somModel.tcam_mask[3][552][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][553][0]=80'h00000000000000c2fbc1;
sos_loop[0].somModel.tcam_mask[3][553][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][554][0]=80'h000000000000004cbb09;
sos_loop[0].somModel.tcam_mask[3][554][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][555][0]=80'h00000000000000ffbbbf;
sos_loop[0].somModel.tcam_mask[3][555][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][556][0]=80'h00000000000000b682c8;
sos_loop[0].somModel.tcam_mask[3][556][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][557][0]=80'h0000000000000052c4da;
sos_loop[0].somModel.tcam_mask[3][557][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][558][0]=80'h00000000000000312a41;
sos_loop[0].somModel.tcam_mask[3][558][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][559][0]=80'h0000000000000008b4d5;
sos_loop[0].somModel.tcam_mask[3][559][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][560][0]=80'h00000000000000f3a2ad;
sos_loop[0].somModel.tcam_mask[3][560][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][561][0]=80'h000000000000006e7c4f;
sos_loop[0].somModel.tcam_mask[3][561][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][562][0]=80'h00000000000000ded8dc;
sos_loop[0].somModel.tcam_mask[3][562][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][563][0]=80'h0000000000000001dc81;
sos_loop[0].somModel.tcam_mask[3][563][0]=80'hfffffffffffffffe0000;
sos_loop[0].somModel.tcam_data[3][564][0]=80'h000000000000000fbaf9;
sos_loop[0].somModel.tcam_mask[3][564][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][565][0]=80'h0000000000000061584b;
sos_loop[0].somModel.tcam_mask[3][565][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][566][0]=80'h000000000000007649b8;
sos_loop[0].somModel.tcam_mask[3][566][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][567][0]=80'h000000000000005f5cd1;
sos_loop[0].somModel.tcam_mask[3][567][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][568][0]=80'h00000000000000f10131;
sos_loop[0].somModel.tcam_mask[3][568][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][569][0]=80'h0000000000000072671c;
sos_loop[0].somModel.tcam_mask[3][569][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][570][0]=80'h00000000000000d3785d;
sos_loop[0].somModel.tcam_mask[3][570][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][571][0]=80'h00000000000000a29593;
sos_loop[0].somModel.tcam_mask[3][571][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][572][0]=80'h00000000000000954c60;
sos_loop[0].somModel.tcam_mask[3][572][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][573][0]=80'h00000000000000c17e8e;
sos_loop[0].somModel.tcam_mask[3][573][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][574][0]=80'h0000000000000009a7ba;
sos_loop[0].somModel.tcam_mask[3][574][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][575][0]=80'h000000000000007072f3;
sos_loop[0].somModel.tcam_mask[3][575][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][576][0]=80'h0000000000000078fcbf;
sos_loop[0].somModel.tcam_mask[3][576][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][577][0]=80'h0000000000000043c1b7;
sos_loop[0].somModel.tcam_mask[3][577][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][578][0]=80'h00000000000000b08007;
sos_loop[0].somModel.tcam_mask[3][578][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][579][0]=80'h00000000000000150566;
sos_loop[0].somModel.tcam_mask[3][579][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][580][0]=80'h00000000000000a9a978;
sos_loop[0].somModel.tcam_mask[3][580][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][581][0]=80'h00000000000000c86b86;
sos_loop[0].somModel.tcam_mask[3][581][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][582][0]=80'h00000000000000f6a9b4;
sos_loop[0].somModel.tcam_mask[3][582][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][583][0]=80'h00000000000000bd5e1d;
sos_loop[0].somModel.tcam_mask[3][583][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][584][0]=80'h000000000000006bdf3d;
sos_loop[0].somModel.tcam_mask[3][584][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][585][0]=80'h000000000000008848ec;
sos_loop[0].somModel.tcam_mask[3][585][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][586][0]=80'h000000000000002de4cb;
sos_loop[0].somModel.tcam_mask[3][586][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][587][0]=80'h00000000000000729081;
sos_loop[0].somModel.tcam_mask[3][587][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][588][0]=80'h000000000000006a8d3d;
sos_loop[0].somModel.tcam_mask[3][588][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][589][0]=80'h00000000000000b986e7;
sos_loop[0].somModel.tcam_mask[3][589][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][590][0]=80'h0000000000000053a9dc;
sos_loop[0].somModel.tcam_mask[3][590][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][591][0]=80'h00000000000000495aab;
sos_loop[0].somModel.tcam_mask[3][591][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][592][0]=80'h000000000000002243c5;
sos_loop[0].somModel.tcam_mask[3][592][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][593][0]=80'h00000000000000932bc5;
sos_loop[0].somModel.tcam_mask[3][593][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][594][0]=80'h00000000000000c7e5a1;
sos_loop[0].somModel.tcam_mask[3][594][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][595][0]=80'h00000000000000519f51;
sos_loop[0].somModel.tcam_mask[3][595][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][596][0]=80'h0000000000000031d9d3;
sos_loop[0].somModel.tcam_mask[3][596][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][597][0]=80'h000000000000006c648c;
sos_loop[0].somModel.tcam_mask[3][597][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][598][0]=80'h00000000000000ca4098;
sos_loop[0].somModel.tcam_mask[3][598][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][599][0]=80'h00000000000000e6aa63;
sos_loop[0].somModel.tcam_mask[3][599][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][600][0]=80'h000000000000009898d6;
sos_loop[0].somModel.tcam_mask[3][600][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][601][0]=80'h000000000000002e0ee6;
sos_loop[0].somModel.tcam_mask[3][601][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][602][0]=80'h000000000000007de959;
sos_loop[0].somModel.tcam_mask[3][602][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][603][0]=80'h0000000000000022ed5e;
sos_loop[0].somModel.tcam_mask[3][603][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][604][0]=80'h00000000000000ef9cd4;
sos_loop[0].somModel.tcam_mask[3][604][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][605][0]=80'h000000000000009e573b;
sos_loop[0].somModel.tcam_mask[3][605][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][606][0]=80'h00000000000000a4a6bf;
sos_loop[0].somModel.tcam_mask[3][606][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][607][0]=80'h0000000000000096fae7;
sos_loop[0].somModel.tcam_mask[3][607][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][608][0]=80'h00000000000000cdbaec;
sos_loop[0].somModel.tcam_mask[3][608][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][609][0]=80'h00000000000000f9a463;
sos_loop[0].somModel.tcam_mask[3][609][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][610][0]=80'h000000000000004e36e0;
sos_loop[0].somModel.tcam_mask[3][610][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][611][0]=80'h00000000000000f0a7a9;
sos_loop[0].somModel.tcam_mask[3][611][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][612][0]=80'h000000000000001ae7e7;
sos_loop[0].somModel.tcam_mask[3][612][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][613][0]=80'h00000000000000facdcc;
sos_loop[0].somModel.tcam_mask[3][613][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][614][0]=80'h00000000000000057f90;
sos_loop[0].somModel.tcam_mask[3][614][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][615][0]=80'h00000000000000b782da;
sos_loop[0].somModel.tcam_mask[3][615][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][616][0]=80'h000000000000000068b3;
sos_loop[0].somModel.tcam_mask[3][616][0]=80'hffffffffffffffff8000;
sos_loop[0].somModel.tcam_data[3][617][0]=80'h000000000000003a8542;
sos_loop[0].somModel.tcam_mask[3][617][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][618][0]=80'h00000000000000662a36;
sos_loop[0].somModel.tcam_mask[3][618][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][619][0]=80'h00000000000000c447e7;
sos_loop[0].somModel.tcam_mask[3][619][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][620][0]=80'h00000000000000428275;
sos_loop[0].somModel.tcam_mask[3][620][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][621][0]=80'h00000000000000207e9f;
sos_loop[0].somModel.tcam_mask[3][621][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][622][0]=80'h00000000000000b5de9b;
sos_loop[0].somModel.tcam_mask[3][622][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][623][0]=80'h00000000000000bdfb18;
sos_loop[0].somModel.tcam_mask[3][623][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][624][0]=80'h000000000000003a7a85;
sos_loop[0].somModel.tcam_mask[3][624][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][625][0]=80'h000000000000006b085d;
sos_loop[0].somModel.tcam_mask[3][625][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][626][0]=80'h00000000000000e56816;
sos_loop[0].somModel.tcam_mask[3][626][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][627][0]=80'h0000000000000018d22b;
sos_loop[0].somModel.tcam_mask[3][627][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][628][0]=80'h00000000000000fd73c1;
sos_loop[0].somModel.tcam_mask[3][628][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][629][0]=80'h00000000000000f65166;
sos_loop[0].somModel.tcam_mask[3][629][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][630][0]=80'h00000000000000aea4f6;
sos_loop[0].somModel.tcam_mask[3][630][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][631][0]=80'h00000000000000378ad7;
sos_loop[0].somModel.tcam_mask[3][631][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][632][0]=80'h000000000000007215cb;
sos_loop[0].somModel.tcam_mask[3][632][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][633][0]=80'h000000000000004370d3;
sos_loop[0].somModel.tcam_mask[3][633][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][634][0]=80'h00000000000000e0bb48;
sos_loop[0].somModel.tcam_mask[3][634][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][635][0]=80'h00000000000000dd2dbc;
sos_loop[0].somModel.tcam_mask[3][635][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][636][0]=80'h00000000000000d10c0d;
sos_loop[0].somModel.tcam_mask[3][636][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][637][0]=80'h0000000000000045ca7b;
sos_loop[0].somModel.tcam_mask[3][637][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][638][0]=80'h0000000000000050ec64;
sos_loop[0].somModel.tcam_mask[3][638][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][639][0]=80'h00000000000000906144;
sos_loop[0].somModel.tcam_mask[3][639][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][640][0]=80'h00000000000000112dc1;
sos_loop[0].somModel.tcam_mask[3][640][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][641][0]=80'h000000000000005b36ae;
sos_loop[0].somModel.tcam_mask[3][641][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][642][0]=80'h000000000000006a5c37;
sos_loop[0].somModel.tcam_mask[3][642][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][643][0]=80'h0000000000000024a942;
sos_loop[0].somModel.tcam_mask[3][643][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][644][0]=80'h00000000000000048e2b;
sos_loop[0].somModel.tcam_mask[3][644][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][645][0]=80'h0000000000000077fa27;
sos_loop[0].somModel.tcam_mask[3][645][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][646][0]=80'h0000000000000078b151;
sos_loop[0].somModel.tcam_mask[3][646][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][647][0]=80'h00000000000000a47604;
sos_loop[0].somModel.tcam_mask[3][647][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][648][0]=80'h00000000000000594a3f;
sos_loop[0].somModel.tcam_mask[3][648][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][649][0]=80'h00000000000000af2e91;
sos_loop[0].somModel.tcam_mask[3][649][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][650][0]=80'h0000000000000054f406;
sos_loop[0].somModel.tcam_mask[3][650][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][651][0]=80'h00000000000000dbd353;
sos_loop[0].somModel.tcam_mask[3][651][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][652][0]=80'h00000000000000a961f7;
sos_loop[0].somModel.tcam_mask[3][652][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][653][0]=80'h00000000000000655384;
sos_loop[0].somModel.tcam_mask[3][653][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][654][0]=80'h0000000000000001b8b2;
sos_loop[0].somModel.tcam_mask[3][654][0]=80'hfffffffffffffffe0000;
sos_loop[0].somModel.tcam_data[3][655][0]=80'h00000000000000b646a0;
sos_loop[0].somModel.tcam_mask[3][655][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][656][0]=80'h00000000000000c35541;
sos_loop[0].somModel.tcam_mask[3][656][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][657][0]=80'h00000000000000aa459d;
sos_loop[0].somModel.tcam_mask[3][657][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][658][0]=80'h00000000000000759b4f;
sos_loop[0].somModel.tcam_mask[3][658][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][659][0]=80'h0000000000000010b764;
sos_loop[0].somModel.tcam_mask[3][659][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][660][0]=80'h000000000000007f2ca2;
sos_loop[0].somModel.tcam_mask[3][660][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][661][0]=80'h00000000000000009605;
sos_loop[0].somModel.tcam_mask[3][661][0]=80'hffffffffffffffff0000;
sos_loop[0].somModel.tcam_data[3][662][0]=80'h00000000000000880ee7;
sos_loop[0].somModel.tcam_mask[3][662][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][663][0]=80'h00000000000000eced99;
sos_loop[0].somModel.tcam_mask[3][663][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][664][0]=80'h000000000000008a05ca;
sos_loop[0].somModel.tcam_mask[3][664][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][665][0]=80'h0000000000000066baf9;
sos_loop[0].somModel.tcam_mask[3][665][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][666][0]=80'h0000000000000096805d;
sos_loop[0].somModel.tcam_mask[3][666][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][667][0]=80'h000000000000000e3de2;
sos_loop[0].somModel.tcam_mask[3][667][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][668][0]=80'h0000000000000015e3df;
sos_loop[0].somModel.tcam_mask[3][668][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][669][0]=80'h00000000000000a47712;
sos_loop[0].somModel.tcam_mask[3][669][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][670][0]=80'h000000000000001932f3;
sos_loop[0].somModel.tcam_mask[3][670][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][671][0]=80'h0000000000000015d54c;
sos_loop[0].somModel.tcam_mask[3][671][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[3][672][0]=80'h000000000000008e6097;
sos_loop[0].somModel.tcam_mask[3][672][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][673][0]=80'h00000000000000026723;
sos_loop[0].somModel.tcam_mask[3][673][0]=80'hfffffffffffffffc0000;
sos_loop[0].somModel.tcam_data[3][674][0]=80'h000000000000002d4201;
sos_loop[0].somModel.tcam_mask[3][674][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][675][0]=80'h0000000000000064a019;
sos_loop[0].somModel.tcam_mask[3][675][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][676][0]=80'h00000000000000052068;
sos_loop[0].somModel.tcam_mask[3][676][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[3][677][0]=80'h000000000000004fc87f;
sos_loop[0].somModel.tcam_mask[3][677][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][678][0]=80'h00000000000000354c4a;
sos_loop[0].somModel.tcam_mask[3][678][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][679][0]=80'h00000000000000c084df;
sos_loop[0].somModel.tcam_mask[3][679][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][680][0]=80'h00000000000000e3af6c;
sos_loop[0].somModel.tcam_mask[3][680][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][681][0]=80'h000000000000009b4c6a;
sos_loop[0].somModel.tcam_mask[3][681][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][682][0]=80'h000000000000004fe061;
sos_loop[0].somModel.tcam_mask[3][682][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][683][0]=80'h00000000000000668b54;
sos_loop[0].somModel.tcam_mask[3][683][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][684][0]=80'h00000000000000b7d2fa;
sos_loop[0].somModel.tcam_mask[3][684][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][685][0]=80'h000000000000007b394b;
sos_loop[0].somModel.tcam_mask[3][685][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][686][0]=80'h00000000000000a0d693;
sos_loop[0].somModel.tcam_mask[3][686][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][687][0]=80'h00000000000000ecb9e8;
sos_loop[0].somModel.tcam_mask[3][687][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][688][0]=80'h00000000000000fa6dcb;
sos_loop[0].somModel.tcam_mask[3][688][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][689][0]=80'h00000000000000549727;
sos_loop[0].somModel.tcam_mask[3][689][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][690][0]=80'h00000000000000563be7;
sos_loop[0].somModel.tcam_mask[3][690][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][691][0]=80'h00000000000000efc0f2;
sos_loop[0].somModel.tcam_mask[3][691][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][692][0]=80'h00000000000000c5e4f2;
sos_loop[0].somModel.tcam_mask[3][692][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][693][0]=80'h0000000000000097e2e2;
sos_loop[0].somModel.tcam_mask[3][693][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][694][0]=80'h00000000000000d71d42;
sos_loop[0].somModel.tcam_mask[3][694][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][695][0]=80'h000000000000002cc08f;
sos_loop[0].somModel.tcam_mask[3][695][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[3][696][0]=80'h000000000000006e18f9;
sos_loop[0].somModel.tcam_mask[3][696][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[3][697][0]=80'h000000000000000fdf59;
sos_loop[0].somModel.tcam_mask[3][697][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[3][698][0]=80'h000000000000008f22b0;
sos_loop[0].somModel.tcam_mask[3][698][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][699][0]=80'h00000000000000f70e50;
sos_loop[0].somModel.tcam_mask[3][699][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[3][700][0]=80'h0000000000000065c364;
sos_loop[0].somModel.tcam_mask[3][700][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.sram_dat[3][0][0]=96'hdeadbf;
sos_loop[0].somModel.sram_ptr[3][0]=939;
sos_loop[0].somModel.sram_dat[3][1][0]=96'hb54f67e3;
sos_loop[0].somModel.sram_ptr[3][1]=3;
sos_loop[0].somModel.sram_dat[3][2][0]=96'h82701ad9;
sos_loop[0].somModel.sram_ptr[3][2]=3;
sos_loop[0].somModel.sram_dat[3][3][0]=96'h73a0f3c7;
sos_loop[0].somModel.sram_ptr[3][3]=3;
sos_loop[0].somModel.sram_dat[3][4][0]=96'h94c7976;
sos_loop[0].somModel.sram_ptr[3][4]=3;
sos_loop[0].somModel.sram_dat[3][5][0]=96'hce105c36;
sos_loop[0].somModel.sram_ptr[3][5]=3;
sos_loop[0].somModel.sram_dat[3][6][0]=96'hb834579a;
sos_loop[0].somModel.sram_ptr[3][6]=3;
sos_loop[0].somModel.sram_dat[3][7][0]=96'h6b75275d;
sos_loop[0].somModel.sram_ptr[3][7]=3;
sos_loop[0].somModel.sram_dat[3][8][0]=96'h65729ff2;
sos_loop[0].somModel.sram_ptr[3][8]=3;
sos_loop[0].somModel.sram_dat[3][9][0]=96'h9c97d69;
sos_loop[0].somModel.sram_ptr[3][9]=3;
sos_loop[0].somModel.sram_dat[3][10][0]=96'h95f0765a;
sos_loop[0].somModel.sram_ptr[3][10]=3;
sos_loop[0].somModel.sram_dat[3][11][0]=96'hc6cb3d40;
sos_loop[0].somModel.sram_ptr[3][11]=3;
sos_loop[0].somModel.sram_dat[3][12][0]=96'h51099d25;
sos_loop[0].somModel.sram_ptr[3][12]=3;
sos_loop[0].somModel.sram_dat[3][13][0]=96'h13be202f;
sos_loop[0].somModel.sram_ptr[3][13]=3;
sos_loop[0].somModel.sram_dat[3][14][0]=96'haded021e;
sos_loop[0].somModel.sram_ptr[3][14]=3;
sos_loop[0].somModel.sram_dat[3][15][0]=96'ha8ab1332;
sos_loop[0].somModel.sram_ptr[3][15]=3;
sos_loop[0].somModel.sram_dat[3][16][0]=96'hdee9be17;
sos_loop[0].somModel.sram_ptr[3][16]=3;
sos_loop[0].somModel.sram_dat[3][17][0]=96'h10344d26;
sos_loop[0].somModel.sram_ptr[3][17]=3;
sos_loop[0].somModel.sram_dat[3][18][0]=96'heee66d45;
sos_loop[0].somModel.sram_ptr[3][18]=3;
sos_loop[0].somModel.sram_dat[3][19][0]=96'h85015a63;
sos_loop[0].somModel.sram_ptr[3][19]=3;
sos_loop[0].somModel.sram_dat[3][20][0]=96'h11b09ad8;
sos_loop[0].somModel.sram_ptr[3][20]=3;
sos_loop[0].somModel.sram_dat[3][21][0]=96'h95ed2ba2;
sos_loop[0].somModel.sram_ptr[3][21]=3;
sos_loop[0].somModel.sram_dat[3][22][0]=96'hae60dfc5;
sos_loop[0].somModel.sram_ptr[3][22]=3;
sos_loop[0].somModel.sram_dat[3][23][0]=96'hf32db0c1;
sos_loop[0].somModel.sram_ptr[3][23]=3;
sos_loop[0].somModel.sram_dat[3][24][0]=96'h9d50520d;
sos_loop[0].somModel.sram_ptr[3][24]=3;
sos_loop[0].somModel.sram_dat[3][25][0]=96'h83fa86a3;
sos_loop[0].somModel.sram_ptr[3][25]=3;
sos_loop[0].somModel.sram_dat[3][26][0]=96'hfed13352;
sos_loop[0].somModel.sram_ptr[3][26]=3;
sos_loop[0].somModel.sram_dat[3][27][0]=96'h6c4cf1a3;
sos_loop[0].somModel.sram_ptr[3][27]=3;
sos_loop[0].somModel.sram_dat[3][28][0]=96'h1e12a2c3;
sos_loop[0].somModel.sram_ptr[3][28]=3;
sos_loop[0].somModel.sram_dat[3][29][0]=96'hb199f9bd;
sos_loop[0].somModel.sram_ptr[3][29]=3;
sos_loop[0].somModel.sram_dat[3][30][0]=96'h5edff01d;
sos_loop[0].somModel.sram_ptr[3][30]=3;
sos_loop[0].somModel.sram_dat[3][31][0]=96'h777705d7;
sos_loop[0].somModel.sram_ptr[3][31]=3;
sos_loop[0].somModel.sram_dat[3][32][0]=96'h65c1fcdf;
sos_loop[0].somModel.sram_ptr[3][32]=3;
sos_loop[0].somModel.sram_dat[3][33][0]=96'h37860217;
sos_loop[0].somModel.sram_ptr[3][33]=3;
sos_loop[0].somModel.sram_dat[3][34][0]=96'h60b3521a;
sos_loop[0].somModel.sram_ptr[3][34]=3;
sos_loop[0].somModel.sram_dat[3][35][0]=96'hd2e417a;
sos_loop[0].somModel.sram_ptr[3][35]=3;
sos_loop[0].somModel.sram_dat[3][36][0]=96'he4f4fa6;
sos_loop[0].somModel.sram_ptr[3][36]=3;
sos_loop[0].somModel.sram_dat[3][37][0]=96'h56ca43a2;
sos_loop[0].somModel.sram_ptr[3][37]=3;
sos_loop[0].somModel.sram_dat[3][38][0]=96'ha3d16cc5;
sos_loop[0].somModel.sram_ptr[3][38]=3;
sos_loop[0].somModel.sram_dat[3][39][0]=96'h17fdfddb;
sos_loop[0].somModel.sram_ptr[3][39]=3;
sos_loop[0].somModel.sram_dat[3][40][0]=96'h8dc5fc1e;
sos_loop[0].somModel.sram_ptr[3][40]=3;
sos_loop[0].somModel.sram_dat[3][41][0]=96'hdda06a7d;
sos_loop[0].somModel.sram_ptr[3][41]=3;
sos_loop[0].somModel.sram_dat[3][42][0]=96'hee1abcfe;
sos_loop[0].somModel.sram_ptr[3][42]=3;
sos_loop[0].somModel.sram_dat[3][43][0]=96'hb6b2c311;
sos_loop[0].somModel.sram_ptr[3][43]=3;
sos_loop[0].somModel.sram_dat[3][44][0]=96'h5222e309;
sos_loop[0].somModel.sram_ptr[3][44]=3;
sos_loop[0].somModel.sram_dat[3][45][0]=96'h4de83400;
sos_loop[0].somModel.sram_ptr[3][45]=3;
sos_loop[0].somModel.sram_dat[3][46][0]=96'hf55ce23a;
sos_loop[0].somModel.sram_ptr[3][46]=3;
sos_loop[0].somModel.sram_dat[3][47][0]=96'h923f30a1;
sos_loop[0].somModel.sram_ptr[3][47]=3;
sos_loop[0].somModel.sram_dat[3][48][0]=96'h2805970;
sos_loop[0].somModel.sram_ptr[3][48]=3;
sos_loop[0].somModel.sram_dat[3][49][0]=96'h600e6cd3;
sos_loop[0].somModel.sram_ptr[3][49]=3;
sos_loop[0].somModel.sram_dat[3][50][0]=96'h560660db;
sos_loop[0].somModel.sram_ptr[3][50]=3;
sos_loop[0].somModel.sram_dat[3][51][0]=96'he78a38a2;
sos_loop[0].somModel.sram_ptr[3][51]=3;
sos_loop[0].somModel.sram_dat[3][52][0]=96'ha2af2509;
sos_loop[0].somModel.sram_ptr[3][52]=3;
sos_loop[0].somModel.sram_dat[3][53][0]=96'hbce83038;
sos_loop[0].somModel.sram_ptr[3][53]=3;
sos_loop[0].somModel.sram_dat[3][54][0]=96'hc6c499c6;
sos_loop[0].somModel.sram_ptr[3][54]=3;
sos_loop[0].somModel.sram_dat[3][55][0]=96'hcfe4fdb8;
sos_loop[0].somModel.sram_ptr[3][55]=3;
sos_loop[0].somModel.sram_dat[3][56][0]=96'he84582e1;
sos_loop[0].somModel.sram_ptr[3][56]=3;
sos_loop[0].somModel.sram_dat[3][57][0]=96'h1cbd8994;
sos_loop[0].somModel.sram_ptr[3][57]=3;
sos_loop[0].somModel.sram_dat[3][58][0]=96'h8725b8fe;
sos_loop[0].somModel.sram_ptr[3][58]=3;
sos_loop[0].somModel.sram_dat[3][59][0]=96'h820f2dae;
sos_loop[0].somModel.sram_ptr[3][59]=3;
sos_loop[0].somModel.sram_dat[3][60][0]=96'hb9ebe16e;
sos_loop[0].somModel.sram_ptr[3][60]=3;
sos_loop[0].somModel.sram_dat[3][61][0]=96'h8f276dcf;
sos_loop[0].somModel.sram_ptr[3][61]=3;
sos_loop[0].somModel.sram_dat[3][62][0]=96'h8158b691;
sos_loop[0].somModel.sram_ptr[3][62]=3;
sos_loop[0].somModel.sram_dat[3][63][0]=96'hf40e5df3;
sos_loop[0].somModel.sram_ptr[3][63]=3;
sos_loop[0].somModel.sram_dat[3][64][0]=96'h7f3fd2ce;
sos_loop[0].somModel.sram_ptr[3][64]=3;
sos_loop[0].somModel.sram_dat[3][65][0]=96'hfb50a4cb;
sos_loop[0].somModel.sram_ptr[3][65]=3;
sos_loop[0].somModel.sram_dat[3][66][0]=96'ha23f290a;
sos_loop[0].somModel.sram_ptr[3][66]=3;
sos_loop[0].somModel.sram_dat[3][67][0]=96'ha249d8fe;
sos_loop[0].somModel.sram_ptr[3][67]=3;
sos_loop[0].somModel.sram_dat[3][68][0]=96'h73ddd4d9;
sos_loop[0].somModel.sram_ptr[3][68]=3;
sos_loop[0].somModel.sram_dat[3][69][0]=96'h3d4518bb;
sos_loop[0].somModel.sram_ptr[3][69]=3;
sos_loop[0].somModel.sram_dat[3][70][0]=96'hb12418a1;
sos_loop[0].somModel.sram_ptr[3][70]=3;
sos_loop[0].somModel.sram_dat[3][71][0]=96'h2b0255f5;
sos_loop[0].somModel.sram_ptr[3][71]=3;
sos_loop[0].somModel.sram_dat[3][72][0]=96'hb26dbe7a;
sos_loop[0].somModel.sram_ptr[3][72]=3;
sos_loop[0].somModel.sram_dat[3][73][0]=96'hbe63e546;
sos_loop[0].somModel.sram_ptr[3][73]=3;
sos_loop[0].somModel.sram_dat[3][74][0]=96'hced8a116;
sos_loop[0].somModel.sram_ptr[3][74]=3;
sos_loop[0].somModel.sram_dat[3][75][0]=96'hd4fd6330;
sos_loop[0].somModel.sram_ptr[3][75]=3;
sos_loop[0].somModel.sram_dat[3][76][0]=96'h89538b5c;
sos_loop[0].somModel.sram_ptr[3][76]=3;
sos_loop[0].somModel.sram_dat[3][77][0]=96'h7545692b;
sos_loop[0].somModel.sram_ptr[3][77]=3;
sos_loop[0].somModel.sram_dat[3][78][0]=96'h6e3d0ccd;
sos_loop[0].somModel.sram_ptr[3][78]=3;
sos_loop[0].somModel.sram_dat[3][79][0]=96'h1f95de86;
sos_loop[0].somModel.sram_ptr[3][79]=3;
sos_loop[0].somModel.sram_dat[3][80][0]=96'h32b5bb45;
sos_loop[0].somModel.sram_ptr[3][80]=3;
sos_loop[0].somModel.sram_dat[3][81][0]=96'hf78ec26e;
sos_loop[0].somModel.sram_ptr[3][81]=3;
sos_loop[0].somModel.sram_dat[3][82][0]=96'h6a4b0fd1;
sos_loop[0].somModel.sram_ptr[3][82]=3;
sos_loop[0].somModel.sram_dat[3][83][0]=96'h1cb2bf20;
sos_loop[0].somModel.sram_ptr[3][83]=3;
sos_loop[0].somModel.sram_dat[3][84][0]=96'hba9bed68;
sos_loop[0].somModel.sram_ptr[3][84]=3;
sos_loop[0].somModel.sram_dat[3][85][0]=96'ha559577e;
sos_loop[0].somModel.sram_ptr[3][85]=3;
sos_loop[0].somModel.sram_dat[3][86][0]=96'h90bad641;
sos_loop[0].somModel.sram_ptr[3][86]=3;
sos_loop[0].somModel.sram_dat[3][87][0]=96'hf6c3245a;
sos_loop[0].somModel.sram_ptr[3][87]=3;
sos_loop[0].somModel.sram_dat[3][88][0]=96'hecda72aa;
sos_loop[0].somModel.sram_ptr[3][88]=3;
sos_loop[0].somModel.sram_dat[3][89][0]=96'hb3b7c2b4;
sos_loop[0].somModel.sram_ptr[3][89]=3;
sos_loop[0].somModel.sram_dat[3][90][0]=96'h1428e333;
sos_loop[0].somModel.sram_ptr[3][90]=3;
sos_loop[0].somModel.sram_dat[3][91][0]=96'h5b902d27;
sos_loop[0].somModel.sram_ptr[3][91]=3;
sos_loop[0].somModel.sram_dat[3][92][0]=96'h153d8c14;
sos_loop[0].somModel.sram_ptr[3][92]=3;
sos_loop[0].somModel.sram_dat[3][93][0]=96'h92d06347;
sos_loop[0].somModel.sram_ptr[3][93]=3;
sos_loop[0].somModel.sram_dat[3][94][0]=96'h2c2c4397;
sos_loop[0].somModel.sram_ptr[3][94]=3;
sos_loop[0].somModel.sram_dat[3][95][0]=96'hb7423e69;
sos_loop[0].somModel.sram_ptr[3][95]=3;
sos_loop[0].somModel.sram_dat[3][96][0]=96'h15a6481;
sos_loop[0].somModel.sram_ptr[3][96]=3;
sos_loop[0].somModel.sram_dat[3][97][0]=96'hdfb988cd;
sos_loop[0].somModel.sram_ptr[3][97]=3;
sos_loop[0].somModel.sram_dat[3][98][0]=96'hcde361c7;
sos_loop[0].somModel.sram_ptr[3][98]=3;
sos_loop[0].somModel.sram_dat[3][99][0]=96'he308f937;
sos_loop[0].somModel.sram_ptr[3][99]=3;
sos_loop[0].somModel.sram_dat[3][100][0]=96'h2164ee50;
sos_loop[0].somModel.sram_ptr[3][100]=3;
sos_loop[0].somModel.sram_dat[3][101][0]=96'h616c5a7f;
sos_loop[0].somModel.sram_ptr[3][101]=3;
sos_loop[0].somModel.sram_dat[3][102][0]=96'hdb1b964e;
sos_loop[0].somModel.sram_ptr[3][102]=3;
sos_loop[0].somModel.sram_dat[3][103][0]=96'h5154a7da;
sos_loop[0].somModel.sram_ptr[3][103]=3;
sos_loop[0].somModel.sram_dat[3][104][0]=96'h5c6ec2c4;
sos_loop[0].somModel.sram_ptr[3][104]=3;
sos_loop[0].somModel.sram_dat[3][105][0]=96'h4294e76d;
sos_loop[0].somModel.sram_ptr[3][105]=3;
sos_loop[0].somModel.sram_dat[3][106][0]=96'h5220f2ca;
sos_loop[0].somModel.sram_ptr[3][106]=3;
sos_loop[0].somModel.sram_dat[3][107][0]=96'hda566993;
sos_loop[0].somModel.sram_ptr[3][107]=3;
sos_loop[0].somModel.sram_dat[3][108][0]=96'h1d318de4;
sos_loop[0].somModel.sram_ptr[3][108]=3;
sos_loop[0].somModel.sram_dat[3][109][0]=96'h3346495f;
sos_loop[0].somModel.sram_ptr[3][109]=3;
sos_loop[0].somModel.sram_dat[3][110][0]=96'hf4a6db31;
sos_loop[0].somModel.sram_ptr[3][110]=3;
sos_loop[0].somModel.sram_dat[3][111][0]=96'h1e9b4645;
sos_loop[0].somModel.sram_ptr[3][111]=3;
sos_loop[0].somModel.sram_dat[3][112][0]=96'hc1ce109e;
sos_loop[0].somModel.sram_ptr[3][112]=3;
sos_loop[0].somModel.sram_dat[3][113][0]=96'h93229de8;
sos_loop[0].somModel.sram_ptr[3][113]=3;
sos_loop[0].somModel.sram_dat[3][114][0]=96'h11553172;
sos_loop[0].somModel.sram_ptr[3][114]=3;
sos_loop[0].somModel.sram_dat[3][115][0]=96'h5db88c38;
sos_loop[0].somModel.sram_ptr[3][115]=3;
sos_loop[0].somModel.sram_dat[3][116][0]=96'h2968364c;
sos_loop[0].somModel.sram_ptr[3][116]=3;
sos_loop[0].somModel.sram_dat[3][117][0]=96'h9c14bafb;
sos_loop[0].somModel.sram_ptr[3][117]=3;
sos_loop[0].somModel.sram_dat[3][118][0]=96'h115ed45f;
sos_loop[0].somModel.sram_ptr[3][118]=3;
sos_loop[0].somModel.sram_dat[3][119][0]=96'hc528fcec;
sos_loop[0].somModel.sram_ptr[3][119]=3;
sos_loop[0].somModel.sram_dat[3][120][0]=96'h2ea562ca;
sos_loop[0].somModel.sram_ptr[3][120]=3;
sos_loop[0].somModel.sram_dat[3][121][0]=96'h70397c26;
sos_loop[0].somModel.sram_ptr[3][121]=3;
sos_loop[0].somModel.sram_dat[3][122][0]=96'h17516503;
sos_loop[0].somModel.sram_ptr[3][122]=3;
sos_loop[0].somModel.sram_dat[3][123][0]=96'he2648a6b;
sos_loop[0].somModel.sram_ptr[3][123]=3;
sos_loop[0].somModel.sram_dat[3][124][0]=96'h9050a552;
sos_loop[0].somModel.sram_ptr[3][124]=3;
sos_loop[0].somModel.sram_dat[3][125][0]=96'h2ae6316d;
sos_loop[0].somModel.sram_ptr[3][125]=3;
sos_loop[0].somModel.sram_dat[3][126][0]=96'h85b27335;
sos_loop[0].somModel.sram_ptr[3][126]=3;
sos_loop[0].somModel.sram_dat[3][127][0]=96'hedcea4e9;
sos_loop[0].somModel.sram_ptr[3][127]=3;
sos_loop[0].somModel.sram_dat[3][128][0]=96'hc3666129;
sos_loop[0].somModel.sram_ptr[3][128]=3;
sos_loop[0].somModel.sram_dat[3][129][0]=96'hdde557c9;
sos_loop[0].somModel.sram_ptr[3][129]=3;
sos_loop[0].somModel.sram_dat[3][130][0]=96'h36fcd376;
sos_loop[0].somModel.sram_ptr[3][130]=3;
sos_loop[0].somModel.sram_dat[3][131][0]=96'hd0642c0d;
sos_loop[0].somModel.sram_ptr[3][131]=3;
sos_loop[0].somModel.sram_dat[3][132][0]=96'h5191ba09;
sos_loop[0].somModel.sram_ptr[3][132]=3;
sos_loop[0].somModel.sram_dat[3][133][0]=96'h307e4946;
sos_loop[0].somModel.sram_ptr[3][133]=3;
sos_loop[0].somModel.sram_dat[3][134][0]=96'h41821824;
sos_loop[0].somModel.sram_ptr[3][134]=3;
sos_loop[0].somModel.sram_dat[3][135][0]=96'h787c80c6;
sos_loop[0].somModel.sram_ptr[3][135]=3;
sos_loop[0].somModel.sram_dat[3][136][0]=96'hf618f71d;
sos_loop[0].somModel.sram_ptr[3][136]=3;
sos_loop[0].somModel.sram_dat[3][137][0]=96'hedacc3d3;
sos_loop[0].somModel.sram_ptr[3][137]=3;
sos_loop[0].somModel.sram_dat[3][138][0]=96'h7e52d942;
sos_loop[0].somModel.sram_ptr[3][138]=3;
sos_loop[0].somModel.sram_dat[3][139][0]=96'h3f71fbaf;
sos_loop[0].somModel.sram_ptr[3][139]=3;
sos_loop[0].somModel.sram_dat[3][140][0]=96'h23350757;
sos_loop[0].somModel.sram_ptr[3][140]=3;
sos_loop[0].somModel.sram_dat[3][141][0]=96'h652439de;
sos_loop[0].somModel.sram_ptr[3][141]=3;
sos_loop[0].somModel.sram_dat[3][142][0]=96'h67c671d1;
sos_loop[0].somModel.sram_ptr[3][142]=3;
sos_loop[0].somModel.sram_dat[3][143][0]=96'h59998fe8;
sos_loop[0].somModel.sram_ptr[3][143]=3;
sos_loop[0].somModel.sram_dat[3][144][0]=96'hd3f88f1f;
sos_loop[0].somModel.sram_ptr[3][144]=3;
sos_loop[0].somModel.sram_dat[3][145][0]=96'hc2b4ab74;
sos_loop[0].somModel.sram_ptr[3][145]=3;
sos_loop[0].somModel.sram_dat[3][146][0]=96'habc85eb1;
sos_loop[0].somModel.sram_ptr[3][146]=3;
sos_loop[0].somModel.sram_dat[3][147][0]=96'h464a1392;
sos_loop[0].somModel.sram_ptr[3][147]=3;
sos_loop[0].somModel.sram_dat[3][148][0]=96'h91c8a041;
sos_loop[0].somModel.sram_ptr[3][148]=3;
sos_loop[0].somModel.sram_dat[3][149][0]=96'h8224a2e1;
sos_loop[0].somModel.sram_ptr[3][149]=3;
sos_loop[0].somModel.sram_dat[3][150][0]=96'he4590888;
sos_loop[0].somModel.sram_ptr[3][150]=3;
sos_loop[0].somModel.sram_dat[3][151][0]=96'hec9ac7c1;
sos_loop[0].somModel.sram_ptr[3][151]=3;
sos_loop[0].somModel.sram_dat[3][152][0]=96'h66424878;
sos_loop[0].somModel.sram_ptr[3][152]=3;
sos_loop[0].somModel.sram_dat[3][153][0]=96'h67af253d;
sos_loop[0].somModel.sram_ptr[3][153]=3;
sos_loop[0].somModel.sram_dat[3][154][0]=96'h45d5dbde;
sos_loop[0].somModel.sram_ptr[3][154]=3;
sos_loop[0].somModel.sram_dat[3][155][0]=96'hc54a488a;
sos_loop[0].somModel.sram_ptr[3][155]=3;
sos_loop[0].somModel.sram_dat[3][156][0]=96'hee973819;
sos_loop[0].somModel.sram_ptr[3][156]=3;
sos_loop[0].somModel.sram_dat[3][157][0]=96'hf58cfd37;
sos_loop[0].somModel.sram_ptr[3][157]=3;
sos_loop[0].somModel.sram_dat[3][158][0]=96'h574bcdc4;
sos_loop[0].somModel.sram_ptr[3][158]=3;
sos_loop[0].somModel.sram_dat[3][159][0]=96'ha7a8595a;
sos_loop[0].somModel.sram_ptr[3][159]=3;
sos_loop[0].somModel.sram_dat[3][160][0]=96'hd3b139e9;
sos_loop[0].somModel.sram_ptr[3][160]=3;
sos_loop[0].somModel.sram_dat[3][161][0]=96'h6e36b346;
sos_loop[0].somModel.sram_ptr[3][161]=3;
sos_loop[0].somModel.sram_dat[3][162][0]=96'hda8acfb4;
sos_loop[0].somModel.sram_ptr[3][162]=3;
sos_loop[0].somModel.sram_dat[3][163][0]=96'h185f3089;
sos_loop[0].somModel.sram_ptr[3][163]=3;
sos_loop[0].somModel.sram_dat[3][164][0]=96'hbde907e3;
sos_loop[0].somModel.sram_ptr[3][164]=3;
sos_loop[0].somModel.sram_dat[3][165][0]=96'h4d5fbad;
sos_loop[0].somModel.sram_ptr[3][165]=3;
sos_loop[0].somModel.sram_dat[3][166][0]=96'hab507ea2;
sos_loop[0].somModel.sram_ptr[3][166]=3;
sos_loop[0].somModel.sram_dat[3][167][0]=96'h6e8feba1;
sos_loop[0].somModel.sram_ptr[3][167]=3;
sos_loop[0].somModel.sram_dat[3][168][0]=96'hd2a5d8f4;
sos_loop[0].somModel.sram_ptr[3][168]=3;
sos_loop[0].somModel.sram_dat[3][169][0]=96'h1f98cf7f;
sos_loop[0].somModel.sram_ptr[3][169]=3;
sos_loop[0].somModel.sram_dat[3][170][0]=96'he00933b5;
sos_loop[0].somModel.sram_ptr[3][170]=3;
sos_loop[0].somModel.sram_dat[3][171][0]=96'h94318208;
sos_loop[0].somModel.sram_ptr[3][171]=3;
sos_loop[0].somModel.sram_dat[3][172][0]=96'h5eef8c5a;
sos_loop[0].somModel.sram_ptr[3][172]=3;
sos_loop[0].somModel.sram_dat[3][173][0]=96'hfb9a2b06;
sos_loop[0].somModel.sram_ptr[3][173]=3;
sos_loop[0].somModel.sram_dat[3][174][0]=96'h1dbc0c13;
sos_loop[0].somModel.sram_ptr[3][174]=3;
sos_loop[0].somModel.sram_dat[3][175][0]=96'h96e2cec1;
sos_loop[0].somModel.sram_ptr[3][175]=3;
sos_loop[0].somModel.sram_dat[3][176][0]=96'hbbfa2397;
sos_loop[0].somModel.sram_ptr[3][176]=3;
sos_loop[0].somModel.sram_dat[3][177][0]=96'h1284be5f;
sos_loop[0].somModel.sram_ptr[3][177]=3;
sos_loop[0].somModel.sram_dat[3][178][0]=96'hb20a2de4;
sos_loop[0].somModel.sram_ptr[3][178]=3;
sos_loop[0].somModel.sram_dat[3][179][0]=96'h521ee751;
sos_loop[0].somModel.sram_ptr[3][179]=3;
sos_loop[0].somModel.sram_dat[3][180][0]=96'h84d1e904;
sos_loop[0].somModel.sram_ptr[3][180]=3;
sos_loop[0].somModel.sram_dat[3][181][0]=96'hbe957768;
sos_loop[0].somModel.sram_ptr[3][181]=3;
sos_loop[0].somModel.sram_dat[3][182][0]=96'h83a7c5dc;
sos_loop[0].somModel.sram_ptr[3][182]=3;
sos_loop[0].somModel.sram_dat[3][183][0]=96'h5ef8ecda;
sos_loop[0].somModel.sram_ptr[3][183]=3;
sos_loop[0].somModel.sram_dat[3][184][0]=96'hc9ef88d4;
sos_loop[0].somModel.sram_ptr[3][184]=3;
sos_loop[0].somModel.sram_dat[3][185][0]=96'hdba7c009;
sos_loop[0].somModel.sram_ptr[3][185]=3;
sos_loop[0].somModel.sram_dat[3][186][0]=96'h6a4242f9;
sos_loop[0].somModel.sram_ptr[3][186]=3;
sos_loop[0].somModel.sram_dat[3][187][0]=96'hcb1f7db1;
sos_loop[0].somModel.sram_ptr[3][187]=3;
sos_loop[0].somModel.sram_dat[3][188][0]=96'h282df15a;
sos_loop[0].somModel.sram_ptr[3][188]=3;
sos_loop[0].somModel.sram_dat[3][189][0]=96'h11da4159;
sos_loop[0].somModel.sram_ptr[3][189]=3;
sos_loop[0].somModel.sram_dat[3][190][0]=96'hc979d2c0;
sos_loop[0].somModel.sram_ptr[3][190]=3;
sos_loop[0].somModel.sram_dat[3][191][0]=96'h15d0a572;
sos_loop[0].somModel.sram_ptr[3][191]=3;
sos_loop[0].somModel.sram_dat[3][192][0]=96'hc90d419a;
sos_loop[0].somModel.sram_ptr[3][192]=3;
sos_loop[0].somModel.sram_dat[3][193][0]=96'hff7786b6;
sos_loop[0].somModel.sram_ptr[3][193]=3;
sos_loop[0].somModel.sram_dat[3][194][0]=96'h694627e0;
sos_loop[0].somModel.sram_ptr[3][194]=3;
sos_loop[0].somModel.sram_dat[3][195][0]=96'h509ecf3e;
sos_loop[0].somModel.sram_ptr[3][195]=3;
sos_loop[0].somModel.sram_dat[3][196][0]=96'h36c22061;
sos_loop[0].somModel.sram_ptr[3][196]=3;
sos_loop[0].somModel.sram_dat[3][197][0]=96'h6df4f696;
sos_loop[0].somModel.sram_ptr[3][197]=3;
sos_loop[0].somModel.sram_dat[3][198][0]=96'h36031f0a;
sos_loop[0].somModel.sram_ptr[3][198]=3;
sos_loop[0].somModel.sram_dat[3][199][0]=96'ha146f76;
sos_loop[0].somModel.sram_ptr[3][199]=3;
sos_loop[0].somModel.sram_dat[3][200][0]=96'hda603da4;
sos_loop[0].somModel.sram_ptr[3][200]=3;
sos_loop[0].somModel.sram_dat[3][201][0]=96'h1bd1cc16;
sos_loop[0].somModel.sram_ptr[3][201]=3;
sos_loop[0].somModel.sram_dat[3][202][0]=96'hb7e843f9;
sos_loop[0].somModel.sram_ptr[3][202]=3;
sos_loop[0].somModel.sram_dat[3][203][0]=96'hba2d6f7;
sos_loop[0].somModel.sram_ptr[3][203]=3;
sos_loop[0].somModel.sram_dat[3][204][0]=96'h51de637b;
sos_loop[0].somModel.sram_ptr[3][204]=3;
sos_loop[0].somModel.sram_dat[3][205][0]=96'h828ec475;
sos_loop[0].somModel.sram_ptr[3][205]=3;
sos_loop[0].somModel.sram_dat[3][206][0]=96'hcf441982;
sos_loop[0].somModel.sram_ptr[3][206]=3;
sos_loop[0].somModel.sram_dat[3][207][0]=96'h6f845ae7;
sos_loop[0].somModel.sram_ptr[3][207]=3;
sos_loop[0].somModel.sram_dat[3][208][0]=96'h86e14992;
sos_loop[0].somModel.sram_ptr[3][208]=3;
sos_loop[0].somModel.sram_dat[3][209][0]=96'hc785a77a;
sos_loop[0].somModel.sram_ptr[3][209]=3;
sos_loop[0].somModel.sram_dat[3][210][0]=96'hf41488dc;
sos_loop[0].somModel.sram_ptr[3][210]=3;
sos_loop[0].somModel.sram_dat[3][211][0]=96'hdc6d7d76;
sos_loop[0].somModel.sram_ptr[3][211]=3;
sos_loop[0].somModel.sram_dat[3][212][0]=96'hb9305c01;
sos_loop[0].somModel.sram_ptr[3][212]=3;
sos_loop[0].somModel.sram_dat[3][213][0]=96'h1b750d7d;
sos_loop[0].somModel.sram_ptr[3][213]=3;
sos_loop[0].somModel.sram_dat[3][214][0]=96'h52e6d13c;
sos_loop[0].somModel.sram_ptr[3][214]=3;
sos_loop[0].somModel.sram_dat[3][215][0]=96'hc8ae7d5e;
sos_loop[0].somModel.sram_ptr[3][215]=3;
sos_loop[0].somModel.sram_dat[3][216][0]=96'hed2db3be;
sos_loop[0].somModel.sram_ptr[3][216]=3;
sos_loop[0].somModel.sram_dat[3][217][0]=96'h66f59500;
sos_loop[0].somModel.sram_ptr[3][217]=3;
sos_loop[0].somModel.sram_dat[3][218][0]=96'h90d448e9;
sos_loop[0].somModel.sram_ptr[3][218]=3;
sos_loop[0].somModel.sram_dat[3][219][0]=96'hb51cbc38;
sos_loop[0].somModel.sram_ptr[3][219]=3;
sos_loop[0].somModel.sram_dat[3][220][0]=96'h47180bae;
sos_loop[0].somModel.sram_ptr[3][220]=3;
sos_loop[0].somModel.sram_dat[3][221][0]=96'he1ffb22b;
sos_loop[0].somModel.sram_ptr[3][221]=3;
sos_loop[0].somModel.sram_dat[3][222][0]=96'heb5391a7;
sos_loop[0].somModel.sram_ptr[3][222]=3;
sos_loop[0].somModel.sram_dat[3][223][0]=96'h1c9a36cd;
sos_loop[0].somModel.sram_ptr[3][223]=3;
sos_loop[0].somModel.sram_dat[3][224][0]=96'h9d48a1ec;
sos_loop[0].somModel.sram_ptr[3][224]=3;
sos_loop[0].somModel.sram_dat[3][225][0]=96'h5163f4bb;
sos_loop[0].somModel.sram_ptr[3][225]=3;
sos_loop[0].somModel.sram_dat[3][226][0]=96'h63169cd6;
sos_loop[0].somModel.sram_ptr[3][226]=3;
sos_loop[0].somModel.sram_dat[3][227][0]=96'hafa075ec;
sos_loop[0].somModel.sram_ptr[3][227]=3;
sos_loop[0].somModel.sram_dat[3][228][0]=96'h100c2296;
sos_loop[0].somModel.sram_ptr[3][228]=3;
sos_loop[0].somModel.sram_dat[3][229][0]=96'hee45cc7a;
sos_loop[0].somModel.sram_ptr[3][229]=3;
sos_loop[0].somModel.sram_dat[3][230][0]=96'h6f92ad29;
sos_loop[0].somModel.sram_ptr[3][230]=3;
sos_loop[0].somModel.sram_dat[3][231][0]=96'h29b9588d;
sos_loop[0].somModel.sram_ptr[3][231]=3;
sos_loop[0].somModel.sram_dat[3][232][0]=96'h618563e7;
sos_loop[0].somModel.sram_ptr[3][232]=3;
sos_loop[0].somModel.sram_dat[3][233][0]=96'ha58cb19c;
sos_loop[0].somModel.sram_ptr[3][233]=3;
sos_loop[0].somModel.sram_dat[3][234][0]=96'h1a5533c0;
sos_loop[0].somModel.sram_ptr[3][234]=3;
sos_loop[0].somModel.sram_dat[3][235][0]=96'h9afdd7cc;
sos_loop[0].somModel.sram_ptr[3][235]=3;
sos_loop[0].somModel.sram_dat[3][236][0]=96'hfb3a8fdc;
sos_loop[0].somModel.sram_ptr[3][236]=3;
sos_loop[0].somModel.sram_dat[3][237][0]=96'h7739a57a;
sos_loop[0].somModel.sram_ptr[3][237]=3;
sos_loop[0].somModel.sram_dat[3][238][0]=96'hbc3079c2;
sos_loop[0].somModel.sram_ptr[3][238]=3;
sos_loop[0].somModel.sram_dat[3][239][0]=96'h566dbe9d;
sos_loop[0].somModel.sram_ptr[3][239]=3;
sos_loop[0].somModel.sram_dat[3][240][0]=96'ha5b90f20;
sos_loop[0].somModel.sram_ptr[3][240]=3;
sos_loop[0].somModel.sram_dat[3][241][0]=96'h17bbd94a;
sos_loop[0].somModel.sram_ptr[3][241]=3;
sos_loop[0].somModel.sram_dat[3][242][0]=96'hd3cf3d16;
sos_loop[0].somModel.sram_ptr[3][242]=3;
sos_loop[0].somModel.sram_dat[3][243][0]=96'h4beeacd4;
sos_loop[0].somModel.sram_ptr[3][243]=3;
sos_loop[0].somModel.sram_dat[3][244][0]=96'h137474a7;
sos_loop[0].somModel.sram_ptr[3][244]=3;
sos_loop[0].somModel.sram_dat[3][245][0]=96'hec022a40;
sos_loop[0].somModel.sram_ptr[3][245]=3;
sos_loop[0].somModel.sram_dat[3][246][0]=96'ha25046c1;
sos_loop[0].somModel.sram_ptr[3][246]=3;
sos_loop[0].somModel.sram_dat[3][247][0]=96'h7035529d;
sos_loop[0].somModel.sram_ptr[3][247]=3;
sos_loop[0].somModel.sram_dat[3][248][0]=96'h1cadbeb4;
sos_loop[0].somModel.sram_ptr[3][248]=3;
sos_loop[0].somModel.sram_dat[3][249][0]=96'h8400df43;
sos_loop[0].somModel.sram_ptr[3][249]=3;
sos_loop[0].somModel.sram_dat[3][250][0]=96'he6b8086f;
sos_loop[0].somModel.sram_ptr[3][250]=3;
sos_loop[0].somModel.sram_dat[3][251][0]=96'h87384f57;
sos_loop[0].somModel.sram_ptr[3][251]=3;
sos_loop[0].somModel.sram_dat[3][252][0]=96'h8d078eb8;
sos_loop[0].somModel.sram_ptr[3][252]=3;
sos_loop[0].somModel.sram_dat[3][253][0]=96'h126db093;
sos_loop[0].somModel.sram_ptr[3][253]=3;
sos_loop[0].somModel.sram_dat[3][254][0]=96'hbf6cb612;
sos_loop[0].somModel.sram_ptr[3][254]=3;
sos_loop[0].somModel.sram_dat[3][255][0]=96'h695c7a60;
sos_loop[0].somModel.sram_ptr[3][255]=3;
sos_loop[0].somModel.sram_dat[3][256][0]=96'h6c8e6262;
sos_loop[0].somModel.sram_ptr[3][256]=3;
sos_loop[0].somModel.sram_dat[3][257][0]=96'h9a4b4a8a;
sos_loop[0].somModel.sram_ptr[3][257]=3;
sos_loop[0].somModel.sram_dat[3][258][0]=96'h9dfaf7d0;
sos_loop[0].somModel.sram_ptr[3][258]=3;
sos_loop[0].somModel.sram_dat[3][259][0]=96'h22388795;
sos_loop[0].somModel.sram_ptr[3][259]=3;
sos_loop[0].somModel.sram_dat[3][260][0]=96'h706887e;
sos_loop[0].somModel.sram_ptr[3][260]=3;
sos_loop[0].somModel.sram_dat[3][261][0]=96'h50674a03;
sos_loop[0].somModel.sram_ptr[3][261]=3;
sos_loop[0].somModel.sram_dat[3][262][0]=96'hc0303373;
sos_loop[0].somModel.sram_ptr[3][262]=3;
sos_loop[0].somModel.sram_dat[3][263][0]=96'h613a337b;
sos_loop[0].somModel.sram_ptr[3][263]=3;
sos_loop[0].somModel.sram_dat[3][264][0]=96'hf56e398f;
sos_loop[0].somModel.sram_ptr[3][264]=3;
sos_loop[0].somModel.sram_dat[3][265][0]=96'h76190ad6;
sos_loop[0].somModel.sram_ptr[3][265]=3;
sos_loop[0].somModel.sram_dat[3][266][0]=96'h1a074b4d;
sos_loop[0].somModel.sram_ptr[3][266]=3;
sos_loop[0].somModel.sram_dat[3][267][0]=96'hb9d382dd;
sos_loop[0].somModel.sram_ptr[3][267]=3;
sos_loop[0].somModel.sram_dat[3][268][0]=96'h49627c77;
sos_loop[0].somModel.sram_ptr[3][268]=3;
sos_loop[0].somModel.sram_dat[3][269][0]=96'h1af7fc78;
sos_loop[0].somModel.sram_ptr[3][269]=3;
sos_loop[0].somModel.sram_dat[3][270][0]=96'h4c5b58c2;
sos_loop[0].somModel.sram_ptr[3][270]=3;
sos_loop[0].somModel.sram_dat[3][271][0]=96'hf7b90362;
sos_loop[0].somModel.sram_ptr[3][271]=3;
sos_loop[0].somModel.sram_dat[3][272][0]=96'h64c19c57;
sos_loop[0].somModel.sram_ptr[3][272]=3;
sos_loop[0].somModel.sram_dat[3][273][0]=96'h4ced0ec5;
sos_loop[0].somModel.sram_ptr[3][273]=3;
sos_loop[0].somModel.sram_dat[3][274][0]=96'h63da1ff4;
sos_loop[0].somModel.sram_ptr[3][274]=3;
sos_loop[0].somModel.sram_dat[3][275][0]=96'hd2bdc987;
sos_loop[0].somModel.sram_ptr[3][275]=3;
sos_loop[0].somModel.sram_dat[3][276][0]=96'h92fa7936;
sos_loop[0].somModel.sram_ptr[3][276]=3;
sos_loop[0].somModel.sram_dat[3][277][0]=96'hf1e9bbdc;
sos_loop[0].somModel.sram_ptr[3][277]=3;
sos_loop[0].somModel.sram_dat[3][278][0]=96'heb9f570f;
sos_loop[0].somModel.sram_ptr[3][278]=3;
sos_loop[0].somModel.sram_dat[3][279][0]=96'h5675f48e;
sos_loop[0].somModel.sram_ptr[3][279]=3;
sos_loop[0].somModel.sram_dat[3][280][0]=96'he73169c;
sos_loop[0].somModel.sram_ptr[3][280]=3;
sos_loop[0].somModel.sram_dat[3][281][0]=96'h12604535;
sos_loop[0].somModel.sram_ptr[3][281]=3;
sos_loop[0].somModel.sram_dat[3][282][0]=96'hf8e3f27b;
sos_loop[0].somModel.sram_ptr[3][282]=3;
sos_loop[0].somModel.sram_dat[3][283][0]=96'h876c9502;
sos_loop[0].somModel.sram_ptr[3][283]=3;
sos_loop[0].somModel.sram_dat[3][284][0]=96'h38ecaf18;
sos_loop[0].somModel.sram_ptr[3][284]=3;
sos_loop[0].somModel.sram_dat[3][285][0]=96'h10bb22bf;
sos_loop[0].somModel.sram_ptr[3][285]=3;
sos_loop[0].somModel.sram_dat[3][286][0]=96'hf4bef27c;
sos_loop[0].somModel.sram_ptr[3][286]=3;
sos_loop[0].somModel.sram_dat[3][287][0]=96'h4cc5a1f3;
sos_loop[0].somModel.sram_ptr[3][287]=3;
sos_loop[0].somModel.sram_dat[3][288][0]=96'hfb03f116;
sos_loop[0].somModel.sram_ptr[3][288]=3;
sos_loop[0].somModel.sram_dat[3][289][0]=96'h1c1d63;
sos_loop[0].somModel.sram_ptr[3][289]=3;
sos_loop[0].somModel.sram_dat[3][290][0]=96'h634ba600;
sos_loop[0].somModel.sram_ptr[3][290]=3;
sos_loop[0].somModel.sram_dat[3][291][0]=96'hb6bfd1ef;
sos_loop[0].somModel.sram_ptr[3][291]=3;
sos_loop[0].somModel.sram_dat[3][292][0]=96'h31a5e63f;
sos_loop[0].somModel.sram_ptr[3][292]=3;
sos_loop[0].somModel.sram_dat[3][293][0]=96'h748ba60c;
sos_loop[0].somModel.sram_ptr[3][293]=3;
sos_loop[0].somModel.sram_dat[3][294][0]=96'h642e6f5e;
sos_loop[0].somModel.sram_ptr[3][294]=3;
sos_loop[0].somModel.sram_dat[3][295][0]=96'h46f2c3d3;
sos_loop[0].somModel.sram_ptr[3][295]=3;
sos_loop[0].somModel.sram_dat[3][296][0]=96'h2636104;
sos_loop[0].somModel.sram_ptr[3][296]=3;
sos_loop[0].somModel.sram_dat[3][297][0]=96'h1ebfe132;
sos_loop[0].somModel.sram_ptr[3][297]=3;
sos_loop[0].somModel.sram_dat[3][298][0]=96'h2b75c41c;
sos_loop[0].somModel.sram_ptr[3][298]=3;
sos_loop[0].somModel.sram_dat[3][299][0]=96'h33c7ddf3;
sos_loop[0].somModel.sram_ptr[3][299]=3;
sos_loop[0].somModel.sram_dat[3][300][0]=96'h9d1dd7c9;
sos_loop[0].somModel.sram_ptr[3][300]=3;
sos_loop[0].somModel.sram_dat[3][301][0]=96'h56c445e5;
sos_loop[0].somModel.sram_ptr[3][301]=3;
sos_loop[0].somModel.sram_dat[3][302][0]=96'h582da58;
sos_loop[0].somModel.sram_ptr[3][302]=3;
sos_loop[0].somModel.sram_dat[3][303][0]=96'h53ea3aa0;
sos_loop[0].somModel.sram_ptr[3][303]=3;
sos_loop[0].somModel.sram_dat[3][304][0]=96'h6528ce42;
sos_loop[0].somModel.sram_ptr[3][304]=3;
sos_loop[0].somModel.sram_dat[3][305][0]=96'ha662e2fd;
sos_loop[0].somModel.sram_ptr[3][305]=3;
sos_loop[0].somModel.sram_dat[3][306][0]=96'h52fcf82a;
sos_loop[0].somModel.sram_ptr[3][306]=3;
sos_loop[0].somModel.sram_dat[3][307][0]=96'ha36b6724;
sos_loop[0].somModel.sram_ptr[3][307]=3;
sos_loop[0].somModel.sram_dat[3][308][0]=96'h57277a34;
sos_loop[0].somModel.sram_ptr[3][308]=3;
sos_loop[0].somModel.sram_dat[3][309][0]=96'h8e243f26;
sos_loop[0].somModel.sram_ptr[3][309]=3;
sos_loop[0].somModel.sram_dat[3][310][0]=96'h3f9a74c6;
sos_loop[0].somModel.sram_ptr[3][310]=3;
sos_loop[0].somModel.sram_dat[3][311][0]=96'h86ae1fea;
sos_loop[0].somModel.sram_ptr[3][311]=3;
sos_loop[0].somModel.sram_dat[3][312][0]=96'h9030da8;
sos_loop[0].somModel.sram_ptr[3][312]=3;
sos_loop[0].somModel.sram_dat[3][313][0]=96'had1f99b7;
sos_loop[0].somModel.sram_ptr[3][313]=3;
sos_loop[0].somModel.sram_dat[3][314][0]=96'h8909580a;
sos_loop[0].somModel.sram_ptr[3][314]=3;
sos_loop[0].somModel.sram_dat[3][315][0]=96'h2ec02701;
sos_loop[0].somModel.sram_ptr[3][315]=3;
sos_loop[0].somModel.sram_dat[3][316][0]=96'h397c1787;
sos_loop[0].somModel.sram_ptr[3][316]=3;
sos_loop[0].somModel.sram_dat[3][317][0]=96'h18384914;
sos_loop[0].somModel.sram_ptr[3][317]=3;
sos_loop[0].somModel.sram_dat[3][318][0]=96'h70844238;
sos_loop[0].somModel.sram_ptr[3][318]=3;
sos_loop[0].somModel.sram_dat[3][319][0]=96'h78d836a6;
sos_loop[0].somModel.sram_ptr[3][319]=3;
sos_loop[0].somModel.sram_dat[3][320][0]=96'h62a813b2;
sos_loop[0].somModel.sram_ptr[3][320]=3;
sos_loop[0].somModel.sram_dat[3][321][0]=96'ha8218af8;
sos_loop[0].somModel.sram_ptr[3][321]=3;
sos_loop[0].somModel.sram_dat[3][322][0]=96'h3fffc90d;
sos_loop[0].somModel.sram_ptr[3][322]=3;
sos_loop[0].somModel.sram_dat[3][323][0]=96'h471270f;
sos_loop[0].somModel.sram_ptr[3][323]=3;
sos_loop[0].somModel.sram_dat[3][324][0]=96'h870c7d6b;
sos_loop[0].somModel.sram_ptr[3][324]=3;
sos_loop[0].somModel.sram_dat[3][325][0]=96'hb1cbd425;
sos_loop[0].somModel.sram_ptr[3][325]=3;
sos_loop[0].somModel.sram_dat[3][326][0]=96'h1ca45b7;
sos_loop[0].somModel.sram_ptr[3][326]=3;
sos_loop[0].somModel.sram_dat[3][327][0]=96'hf9b10ce0;
sos_loop[0].somModel.sram_ptr[3][327]=3;
sos_loop[0].somModel.sram_dat[3][328][0]=96'h5bc3d7cc;
sos_loop[0].somModel.sram_ptr[3][328]=3;
sos_loop[0].somModel.sram_dat[3][329][0]=96'h78b9b3f0;
sos_loop[0].somModel.sram_ptr[3][329]=3;
sos_loop[0].somModel.sram_dat[3][330][0]=96'hd4aa27c8;
sos_loop[0].somModel.sram_ptr[3][330]=3;
sos_loop[0].somModel.sram_dat[3][331][0]=96'h5f341aa9;
sos_loop[0].somModel.sram_ptr[3][331]=3;
sos_loop[0].somModel.sram_dat[3][332][0]=96'hba354357;
sos_loop[0].somModel.sram_ptr[3][332]=3;
sos_loop[0].somModel.sram_dat[3][333][0]=96'h88c143b0;
sos_loop[0].somModel.sram_ptr[3][333]=3;
sos_loop[0].somModel.sram_dat[3][334][0]=96'h48d9a0b4;
sos_loop[0].somModel.sram_ptr[3][334]=3;
sos_loop[0].somModel.sram_dat[3][335][0]=96'hab4daf75;
sos_loop[0].somModel.sram_ptr[3][335]=3;
sos_loop[0].somModel.sram_dat[3][336][0]=96'hd975a916;
sos_loop[0].somModel.sram_ptr[3][336]=3;
sos_loop[0].somModel.sram_dat[3][337][0]=96'he845c902;
sos_loop[0].somModel.sram_ptr[3][337]=3;
sos_loop[0].somModel.sram_dat[3][338][0]=96'h878c2f86;
sos_loop[0].somModel.sram_ptr[3][338]=3;
sos_loop[0].somModel.sram_dat[3][339][0]=96'hba02f376;
sos_loop[0].somModel.sram_ptr[3][339]=3;
sos_loop[0].somModel.sram_dat[3][340][0]=96'hfe0f25ec;
sos_loop[0].somModel.sram_ptr[3][340]=3;
sos_loop[0].somModel.sram_dat[3][341][0]=96'hbcce8db5;
sos_loop[0].somModel.sram_ptr[3][341]=3;
sos_loop[0].somModel.sram_dat[3][342][0]=96'hc3cb15c5;
sos_loop[0].somModel.sram_ptr[3][342]=3;
sos_loop[0].somModel.sram_dat[3][343][0]=96'h32042660;
sos_loop[0].somModel.sram_ptr[3][343]=3;
sos_loop[0].somModel.sram_dat[3][344][0]=96'h713fad01;
sos_loop[0].somModel.sram_ptr[3][344]=3;
sos_loop[0].somModel.sram_dat[3][345][0]=96'h1e45babb;
sos_loop[0].somModel.sram_ptr[3][345]=3;
sos_loop[0].somModel.sram_dat[3][346][0]=96'h537ea7b5;
sos_loop[0].somModel.sram_ptr[3][346]=3;
sos_loop[0].somModel.sram_dat[3][347][0]=96'h2451b99d;
sos_loop[0].somModel.sram_ptr[3][347]=3;
sos_loop[0].somModel.sram_dat[3][348][0]=96'h8c16bba1;
sos_loop[0].somModel.sram_ptr[3][348]=3;
sos_loop[0].somModel.sram_dat[3][349][0]=96'ha6d92913;
sos_loop[0].somModel.sram_ptr[3][349]=3;
sos_loop[0].somModel.sram_dat[3][350][0]=96'hc44e2eee;
sos_loop[0].somModel.sram_ptr[3][350]=3;
sos_loop[0].somModel.sram_dat[3][351][0]=96'h9f76d085;
sos_loop[0].somModel.sram_ptr[3][351]=3;
sos_loop[0].somModel.sram_dat[3][352][0]=96'h774bd3b;
sos_loop[0].somModel.sram_ptr[3][352]=3;
sos_loop[0].somModel.sram_dat[3][353][0]=96'hb8c9750b;
sos_loop[0].somModel.sram_ptr[3][353]=3;
sos_loop[0].somModel.sram_dat[3][354][0]=96'h3b9ced0c;
sos_loop[0].somModel.sram_ptr[3][354]=3;
sos_loop[0].somModel.sram_dat[3][355][0]=96'he822c48d;
sos_loop[0].somModel.sram_ptr[3][355]=3;
sos_loop[0].somModel.sram_dat[3][356][0]=96'h605c12f0;
sos_loop[0].somModel.sram_ptr[3][356]=3;
sos_loop[0].somModel.sram_dat[3][357][0]=96'hd1c12819;
sos_loop[0].somModel.sram_ptr[3][357]=3;
sos_loop[0].somModel.sram_dat[3][358][0]=96'h48d1d320;
sos_loop[0].somModel.sram_ptr[3][358]=3;
sos_loop[0].somModel.sram_dat[3][359][0]=96'h3b2aa084;
sos_loop[0].somModel.sram_ptr[3][359]=3;
sos_loop[0].somModel.sram_dat[3][360][0]=96'h16bb4af9;
sos_loop[0].somModel.sram_ptr[3][360]=3;
sos_loop[0].somModel.sram_dat[3][361][0]=96'hfab919eb;
sos_loop[0].somModel.sram_ptr[3][361]=3;
sos_loop[0].somModel.sram_dat[3][362][0]=96'h9632817;
sos_loop[0].somModel.sram_ptr[3][362]=3;
sos_loop[0].somModel.sram_dat[3][363][0]=96'h2a14c3c5;
sos_loop[0].somModel.sram_ptr[3][363]=3;
sos_loop[0].somModel.sram_dat[3][364][0]=96'h88430aa;
sos_loop[0].somModel.sram_ptr[3][364]=3;
sos_loop[0].somModel.sram_dat[3][365][0]=96'h4b138290;
sos_loop[0].somModel.sram_ptr[3][365]=3;
sos_loop[0].somModel.sram_dat[3][366][0]=96'ha4328192;
sos_loop[0].somModel.sram_ptr[3][366]=3;
sos_loop[0].somModel.sram_dat[3][367][0]=96'haf74e5f0;
sos_loop[0].somModel.sram_ptr[3][367]=3;
sos_loop[0].somModel.sram_dat[3][368][0]=96'hadcbcea6;
sos_loop[0].somModel.sram_ptr[3][368]=3;
sos_loop[0].somModel.sram_dat[3][369][0]=96'h95e27aa3;
sos_loop[0].somModel.sram_ptr[3][369]=3;
sos_loop[0].somModel.sram_dat[3][370][0]=96'h2f201bf5;
sos_loop[0].somModel.sram_ptr[3][370]=3;
sos_loop[0].somModel.sram_dat[3][371][0]=96'ha17dce45;
sos_loop[0].somModel.sram_ptr[3][371]=3;
sos_loop[0].somModel.sram_dat[3][372][0]=96'h9267213c;
sos_loop[0].somModel.sram_ptr[3][372]=3;
sos_loop[0].somModel.sram_dat[3][373][0]=96'h2307fd2f;
sos_loop[0].somModel.sram_ptr[3][373]=3;
sos_loop[0].somModel.sram_dat[3][374][0]=96'hf7c0c8ec;
sos_loop[0].somModel.sram_ptr[3][374]=3;
sos_loop[0].somModel.sram_dat[3][375][0]=96'hc01c6536;
sos_loop[0].somModel.sram_ptr[3][375]=3;
sos_loop[0].somModel.sram_dat[3][376][0]=96'h5821ab3b;
sos_loop[0].somModel.sram_ptr[3][376]=3;
sos_loop[0].somModel.sram_dat[3][377][0]=96'h393a4f1e;
sos_loop[0].somModel.sram_ptr[3][377]=3;
sos_loop[0].somModel.sram_dat[3][378][0]=96'h4ccacbaa;
sos_loop[0].somModel.sram_ptr[3][378]=3;
sos_loop[0].somModel.sram_dat[3][379][0]=96'hbb0cce2;
sos_loop[0].somModel.sram_ptr[3][379]=3;
sos_loop[0].somModel.sram_dat[3][380][0]=96'h4a3557dc;
sos_loop[0].somModel.sram_ptr[3][380]=3;
sos_loop[0].somModel.sram_dat[3][381][0]=96'ha7f5f126;
sos_loop[0].somModel.sram_ptr[3][381]=3;
sos_loop[0].somModel.sram_dat[3][382][0]=96'hecbf5817;
sos_loop[0].somModel.sram_ptr[3][382]=3;
sos_loop[0].somModel.sram_dat[3][383][0]=96'h4fcce4ae;
sos_loop[0].somModel.sram_ptr[3][383]=3;
sos_loop[0].somModel.sram_dat[3][384][0]=96'h49ca82c1;
sos_loop[0].somModel.sram_ptr[3][384]=3;
sos_loop[0].somModel.sram_dat[3][385][0]=96'hc256a85f;
sos_loop[0].somModel.sram_ptr[3][385]=3;
sos_loop[0].somModel.sram_dat[3][386][0]=96'hd0e74b83;
sos_loop[0].somModel.sram_ptr[3][386]=3;
sos_loop[0].somModel.sram_dat[3][387][0]=96'hf790724d;
sos_loop[0].somModel.sram_ptr[3][387]=3;
sos_loop[0].somModel.sram_dat[3][388][0]=96'haa4fdd5a;
sos_loop[0].somModel.sram_ptr[3][388]=3;
sos_loop[0].somModel.sram_dat[3][389][0]=96'h9302e606;
sos_loop[0].somModel.sram_ptr[3][389]=3;
sos_loop[0].somModel.sram_dat[3][390][0]=96'h774c0a95;
sos_loop[0].somModel.sram_ptr[3][390]=3;
sos_loop[0].somModel.sram_dat[3][391][0]=96'hfe7ba7a6;
sos_loop[0].somModel.sram_ptr[3][391]=3;
sos_loop[0].somModel.sram_dat[3][392][0]=96'h763c92c9;
sos_loop[0].somModel.sram_ptr[3][392]=3;
sos_loop[0].somModel.sram_dat[3][393][0]=96'h161007b1;
sos_loop[0].somModel.sram_ptr[3][393]=3;
sos_loop[0].somModel.sram_dat[3][394][0]=96'h2a09f69b;
sos_loop[0].somModel.sram_ptr[3][394]=3;
sos_loop[0].somModel.sram_dat[3][395][0]=96'h8f0631a;
sos_loop[0].somModel.sram_ptr[3][395]=3;
sos_loop[0].somModel.sram_dat[3][396][0]=96'h6e5a5a64;
sos_loop[0].somModel.sram_ptr[3][396]=3;
sos_loop[0].somModel.sram_dat[3][397][0]=96'he4f1fdf8;
sos_loop[0].somModel.sram_ptr[3][397]=3;
sos_loop[0].somModel.sram_dat[3][398][0]=96'h82ee13b8;
sos_loop[0].somModel.sram_ptr[3][398]=3;
sos_loop[0].somModel.sram_dat[3][399][0]=96'h3ebac666;
sos_loop[0].somModel.sram_ptr[3][399]=3;
sos_loop[0].somModel.sram_dat[3][400][0]=96'hc30bb880;
sos_loop[0].somModel.sram_ptr[3][400]=3;
sos_loop[0].somModel.sram_dat[3][401][0]=96'h7bd0807a;
sos_loop[0].somModel.sram_ptr[3][401]=3;
sos_loop[0].somModel.sram_dat[3][402][0]=96'h69c9a36a;
sos_loop[0].somModel.sram_ptr[3][402]=3;
sos_loop[0].somModel.sram_dat[3][403][0]=96'h6dfa7ea1;
sos_loop[0].somModel.sram_ptr[3][403]=3;
sos_loop[0].somModel.sram_dat[3][404][0]=96'h465e2174;
sos_loop[0].somModel.sram_ptr[3][404]=3;
sos_loop[0].somModel.sram_dat[3][405][0]=96'hd690c48f;
sos_loop[0].somModel.sram_ptr[3][405]=3;
sos_loop[0].somModel.sram_dat[3][406][0]=96'h4dfb8bb3;
sos_loop[0].somModel.sram_ptr[3][406]=3;
sos_loop[0].somModel.sram_dat[3][407][0]=96'hfcfb8a1d;
sos_loop[0].somModel.sram_ptr[3][407]=3;
sos_loop[0].somModel.sram_dat[3][408][0]=96'h1e97dfa7;
sos_loop[0].somModel.sram_ptr[3][408]=3;
sos_loop[0].somModel.sram_dat[3][409][0]=96'hfb45ee29;
sos_loop[0].somModel.sram_ptr[3][409]=3;
sos_loop[0].somModel.sram_dat[3][410][0]=96'h2e75bd78;
sos_loop[0].somModel.sram_ptr[3][410]=3;
sos_loop[0].somModel.sram_dat[3][411][0]=96'h22c82a03;
sos_loop[0].somModel.sram_ptr[3][411]=3;
sos_loop[0].somModel.sram_dat[3][412][0]=96'hb5e57ae6;
sos_loop[0].somModel.sram_ptr[3][412]=3;
sos_loop[0].somModel.sram_dat[3][413][0]=96'h6d61818d;
sos_loop[0].somModel.sram_ptr[3][413]=3;
sos_loop[0].somModel.sram_dat[3][414][0]=96'h89bd817f;
sos_loop[0].somModel.sram_ptr[3][414]=3;
sos_loop[0].somModel.sram_dat[3][415][0]=96'h39a3e363;
sos_loop[0].somModel.sram_ptr[3][415]=3;
sos_loop[0].somModel.sram_dat[3][416][0]=96'hf1d02dcb;
sos_loop[0].somModel.sram_ptr[3][416]=3;
sos_loop[0].somModel.sram_dat[3][417][0]=96'he7cab4e5;
sos_loop[0].somModel.sram_ptr[3][417]=3;
sos_loop[0].somModel.sram_dat[3][418][0]=96'h93c91bc5;
sos_loop[0].somModel.sram_ptr[3][418]=3;
sos_loop[0].somModel.sram_dat[3][419][0]=96'h7e18e057;
sos_loop[0].somModel.sram_ptr[3][419]=3;
sos_loop[0].somModel.sram_dat[3][420][0]=96'ha32ff2f6;
sos_loop[0].somModel.sram_ptr[3][420]=3;
sos_loop[0].somModel.sram_dat[3][421][0]=96'h176b62ce;
sos_loop[0].somModel.sram_ptr[3][421]=3;
sos_loop[0].somModel.sram_dat[3][422][0]=96'h31482dc2;
sos_loop[0].somModel.sram_ptr[3][422]=3;
sos_loop[0].somModel.sram_dat[3][423][0]=96'h5dd0192c;
sos_loop[0].somModel.sram_ptr[3][423]=3;
sos_loop[0].somModel.sram_dat[3][424][0]=96'h9c37fed2;
sos_loop[0].somModel.sram_ptr[3][424]=3;
sos_loop[0].somModel.sram_dat[3][425][0]=96'h4172ae7a;
sos_loop[0].somModel.sram_ptr[3][425]=3;
sos_loop[0].somModel.sram_dat[3][426][0]=96'h7a4b700b;
sos_loop[0].somModel.sram_ptr[3][426]=3;
sos_loop[0].somModel.sram_dat[3][427][0]=96'h5b6bae30;
sos_loop[0].somModel.sram_ptr[3][427]=3;
sos_loop[0].somModel.sram_dat[3][428][0]=96'hc829489d;
sos_loop[0].somModel.sram_ptr[3][428]=3;
sos_loop[0].somModel.sram_dat[3][429][0]=96'h1fe9c4aa;
sos_loop[0].somModel.sram_ptr[3][429]=3;
sos_loop[0].somModel.sram_dat[3][430][0]=96'h455925b1;
sos_loop[0].somModel.sram_ptr[3][430]=3;
sos_loop[0].somModel.sram_dat[3][431][0]=96'heec3172f;
sos_loop[0].somModel.sram_ptr[3][431]=3;
sos_loop[0].somModel.sram_dat[3][432][0]=96'hbe5b95ba;
sos_loop[0].somModel.sram_ptr[3][432]=3;
sos_loop[0].somModel.sram_dat[3][433][0]=96'hf7c5318d;
sos_loop[0].somModel.sram_ptr[3][433]=3;
sos_loop[0].somModel.sram_dat[3][434][0]=96'h32b3ab3d;
sos_loop[0].somModel.sram_ptr[3][434]=3;
sos_loop[0].somModel.sram_dat[3][435][0]=96'hf03288ba;
sos_loop[0].somModel.sram_ptr[3][435]=3;
sos_loop[0].somModel.sram_dat[3][436][0]=96'h54d26dab;
sos_loop[0].somModel.sram_ptr[3][436]=3;
sos_loop[0].somModel.sram_dat[3][437][0]=96'h3b35ba0b;
sos_loop[0].somModel.sram_ptr[3][437]=3;
sos_loop[0].somModel.sram_dat[3][438][0]=96'h4725d7df;
sos_loop[0].somModel.sram_ptr[3][438]=3;
sos_loop[0].somModel.sram_dat[3][439][0]=96'h82bd2740;
sos_loop[0].somModel.sram_ptr[3][439]=3;
sos_loop[0].somModel.sram_dat[3][440][0]=96'h4ab16fe6;
sos_loop[0].somModel.sram_ptr[3][440]=3;
sos_loop[0].somModel.sram_dat[3][441][0]=96'hb8828761;
sos_loop[0].somModel.sram_ptr[3][441]=3;
sos_loop[0].somModel.sram_dat[3][442][0]=96'hd7fed41e;
sos_loop[0].somModel.sram_ptr[3][442]=3;
sos_loop[0].somModel.sram_dat[3][443][0]=96'h927e89c8;
sos_loop[0].somModel.sram_ptr[3][443]=3;
sos_loop[0].somModel.sram_dat[3][444][0]=96'h69ce648c;
sos_loop[0].somModel.sram_ptr[3][444]=3;
sos_loop[0].somModel.sram_dat[3][445][0]=96'ha98af6be;
sos_loop[0].somModel.sram_ptr[3][445]=3;
sos_loop[0].somModel.sram_dat[3][446][0]=96'h830c2297;
sos_loop[0].somModel.sram_ptr[3][446]=3;
sos_loop[0].somModel.sram_dat[3][447][0]=96'h8a7c096a;
sos_loop[0].somModel.sram_ptr[3][447]=3;
sos_loop[0].somModel.sram_dat[3][448][0]=96'h87b80521;
sos_loop[0].somModel.sram_ptr[3][448]=3;
sos_loop[0].somModel.sram_dat[3][449][0]=96'h7b3a4eaa;
sos_loop[0].somModel.sram_ptr[3][449]=3;
sos_loop[0].somModel.sram_dat[3][450][0]=96'hbe3050db;
sos_loop[0].somModel.sram_ptr[3][450]=3;
sos_loop[0].somModel.sram_dat[3][451][0]=96'hdc28e522;
sos_loop[0].somModel.sram_ptr[3][451]=3;
sos_loop[0].somModel.sram_dat[3][452][0]=96'h36b04f1c;
sos_loop[0].somModel.sram_ptr[3][452]=3;
sos_loop[0].somModel.sram_dat[3][453][0]=96'h403a7c3e;
sos_loop[0].somModel.sram_ptr[3][453]=3;
sos_loop[0].somModel.sram_dat[3][454][0]=96'h3955090;
sos_loop[0].somModel.sram_ptr[3][454]=3;
sos_loop[0].somModel.sram_dat[3][455][0]=96'h9b0e15b;
sos_loop[0].somModel.sram_ptr[3][455]=3;
sos_loop[0].somModel.sram_dat[3][456][0]=96'h9d7eb941;
sos_loop[0].somModel.sram_ptr[3][456]=3;
sos_loop[0].somModel.sram_dat[3][457][0]=96'h92cc7b97;
sos_loop[0].somModel.sram_ptr[3][457]=3;
sos_loop[0].somModel.sram_dat[3][458][0]=96'h526e091b;
sos_loop[0].somModel.sram_ptr[3][458]=3;
sos_loop[0].somModel.sram_dat[3][459][0]=96'h3f5d769e;
sos_loop[0].somModel.sram_ptr[3][459]=3;
sos_loop[0].somModel.sram_dat[3][460][0]=96'h150c92e2;
sos_loop[0].somModel.sram_ptr[3][460]=3;
sos_loop[0].somModel.sram_dat[3][461][0]=96'he834138a;
sos_loop[0].somModel.sram_ptr[3][461]=3;
sos_loop[0].somModel.sram_dat[3][462][0]=96'hc34ca9d1;
sos_loop[0].somModel.sram_ptr[3][462]=3;
sos_loop[0].somModel.sram_dat[3][463][0]=96'hb3572efe;
sos_loop[0].somModel.sram_ptr[3][463]=3;
sos_loop[0].somModel.sram_dat[3][464][0]=96'hc6f229f9;
sos_loop[0].somModel.sram_ptr[3][464]=3;
sos_loop[0].somModel.sram_dat[3][465][0]=96'he5cbabe9;
sos_loop[0].somModel.sram_ptr[3][465]=3;
sos_loop[0].somModel.sram_dat[3][466][0]=96'h864f25f7;
sos_loop[0].somModel.sram_ptr[3][466]=3;
sos_loop[0].somModel.sram_dat[3][467][0]=96'h67c4066d;
sos_loop[0].somModel.sram_ptr[3][467]=3;
sos_loop[0].somModel.sram_dat[3][468][0]=96'h9de1cb00;
sos_loop[0].somModel.sram_ptr[3][468]=3;
sos_loop[0].somModel.sram_dat[3][469][0]=96'h34248c05;
sos_loop[0].somModel.sram_ptr[3][469]=3;
sos_loop[0].somModel.sram_dat[3][470][0]=96'hc58b25e4;
sos_loop[0].somModel.sram_ptr[3][470]=3;
sos_loop[0].somModel.sram_dat[3][471][0]=96'hb3f968f6;
sos_loop[0].somModel.sram_ptr[3][471]=3;
sos_loop[0].somModel.sram_dat[3][472][0]=96'h8948dfa0;
sos_loop[0].somModel.sram_ptr[3][472]=3;
sos_loop[0].somModel.sram_dat[3][473][0]=96'h6186b4d5;
sos_loop[0].somModel.sram_ptr[3][473]=3;
sos_loop[0].somModel.sram_dat[3][474][0]=96'he5423ca6;
sos_loop[0].somModel.sram_ptr[3][474]=3;
sos_loop[0].somModel.sram_dat[3][475][0]=96'hfb755c87;
sos_loop[0].somModel.sram_ptr[3][475]=3;
sos_loop[0].somModel.sram_dat[3][476][0]=96'ha2792929;
sos_loop[0].somModel.sram_ptr[3][476]=3;
sos_loop[0].somModel.sram_dat[3][477][0]=96'hd4bca2bb;
sos_loop[0].somModel.sram_ptr[3][477]=3;
sos_loop[0].somModel.sram_dat[3][478][0]=96'h3c15896e;
sos_loop[0].somModel.sram_ptr[3][478]=3;
sos_loop[0].somModel.sram_dat[3][479][0]=96'h88e915d3;
sos_loop[0].somModel.sram_ptr[3][479]=3;
sos_loop[0].somModel.sram_dat[3][480][0]=96'h62db80d6;
sos_loop[0].somModel.sram_ptr[3][480]=3;
sos_loop[0].somModel.sram_dat[3][481][0]=96'h4c481bbc;
sos_loop[0].somModel.sram_ptr[3][481]=3;
sos_loop[0].somModel.sram_dat[3][482][0]=96'h9dbbbd6;
sos_loop[0].somModel.sram_ptr[3][482]=3;
sos_loop[0].somModel.sram_dat[3][483][0]=96'hfcce66eb;
sos_loop[0].somModel.sram_ptr[3][483]=3;
sos_loop[0].somModel.sram_dat[3][484][0]=96'h6830b811;
sos_loop[0].somModel.sram_ptr[3][484]=3;
sos_loop[0].somModel.sram_dat[3][485][0]=96'h4379b461;
sos_loop[0].somModel.sram_ptr[3][485]=3;
sos_loop[0].somModel.sram_dat[3][486][0]=96'h68938af3;
sos_loop[0].somModel.sram_ptr[3][486]=3;
sos_loop[0].somModel.sram_dat[3][487][0]=96'h7ff6250d;
sos_loop[0].somModel.sram_ptr[3][487]=3;
sos_loop[0].somModel.sram_dat[3][488][0]=96'hd0b2e426;
sos_loop[0].somModel.sram_ptr[3][488]=3;
sos_loop[0].somModel.sram_dat[3][489][0]=96'he0769eb3;
sos_loop[0].somModel.sram_ptr[3][489]=3;
sos_loop[0].somModel.sram_dat[3][490][0]=96'hebca488e;
sos_loop[0].somModel.sram_ptr[3][490]=3;
sos_loop[0].somModel.sram_dat[3][491][0]=96'ha7d59609;
sos_loop[0].somModel.sram_ptr[3][491]=3;
sos_loop[0].somModel.sram_dat[3][492][0]=96'h861d983b;
sos_loop[0].somModel.sram_ptr[3][492]=3;
sos_loop[0].somModel.sram_dat[3][493][0]=96'h13c0f8ae;
sos_loop[0].somModel.sram_ptr[3][493]=3;
sos_loop[0].somModel.sram_dat[3][494][0]=96'h9aac6fda;
sos_loop[0].somModel.sram_ptr[3][494]=3;
sos_loop[0].somModel.sram_dat[3][495][0]=96'h43d9df1c;
sos_loop[0].somModel.sram_ptr[3][495]=3;
sos_loop[0].somModel.sram_dat[3][496][0]=96'he9a06c24;
sos_loop[0].somModel.sram_ptr[3][496]=3;
sos_loop[0].somModel.sram_dat[3][497][0]=96'hac0241b2;
sos_loop[0].somModel.sram_ptr[3][497]=3;
sos_loop[0].somModel.sram_dat[3][498][0]=96'h7612253b;
sos_loop[0].somModel.sram_ptr[3][498]=3;
sos_loop[0].somModel.sram_dat[3][499][0]=96'hed8abb5c;
sos_loop[0].somModel.sram_ptr[3][499]=3;
sos_loop[0].somModel.sram_dat[3][500][0]=96'h6f9d5e51;
sos_loop[0].somModel.sram_ptr[3][500]=3;
sos_loop[0].somModel.sram_dat[3][501][0]=96'h16ac4efe;
sos_loop[0].somModel.sram_ptr[3][501]=3;
sos_loop[0].somModel.sram_dat[3][502][0]=96'hc3ab0255;
sos_loop[0].somModel.sram_ptr[3][502]=3;
sos_loop[0].somModel.sram_dat[3][503][0]=96'hc4f30409;
sos_loop[0].somModel.sram_ptr[3][503]=3;
sos_loop[0].somModel.sram_dat[3][504][0]=96'h39a47d32;
sos_loop[0].somModel.sram_ptr[3][504]=3;
sos_loop[0].somModel.sram_dat[3][505][0]=96'h935c5f96;
sos_loop[0].somModel.sram_ptr[3][505]=3;
sos_loop[0].somModel.sram_dat[3][506][0]=96'h46b4c54a;
sos_loop[0].somModel.sram_ptr[3][506]=3;
sos_loop[0].somModel.sram_dat[3][507][0]=96'h94b72783;
sos_loop[0].somModel.sram_ptr[3][507]=3;
sos_loop[0].somModel.sram_dat[3][508][0]=96'hb1299113;
sos_loop[0].somModel.sram_ptr[3][508]=3;
sos_loop[0].somModel.sram_dat[3][509][0]=96'h8bed837b;
sos_loop[0].somModel.sram_ptr[3][509]=3;
sos_loop[0].somModel.sram_dat[3][510][0]=96'h4420d131;
sos_loop[0].somModel.sram_ptr[3][510]=3;
sos_loop[0].somModel.sram_dat[3][511][0]=96'h53eb678a;
sos_loop[0].somModel.sram_ptr[3][511]=3;
sos_loop[0].somModel.sram_dat[3][512][0]=96'hbae75dd5;
sos_loop[0].somModel.sram_ptr[3][512]=3;
sos_loop[0].somModel.sram_dat[3][513][0]=96'h18f29af4;
sos_loop[0].somModel.sram_ptr[3][513]=3;
sos_loop[0].somModel.sram_dat[3][514][0]=96'h34bf20e6;
sos_loop[0].somModel.sram_ptr[3][514]=3;
sos_loop[0].somModel.sram_dat[3][515][0]=96'hd7e1bf9e;
sos_loop[0].somModel.sram_ptr[3][515]=3;
sos_loop[0].somModel.sram_dat[3][516][0]=96'hc653b4a2;
sos_loop[0].somModel.sram_ptr[3][516]=3;
sos_loop[0].somModel.sram_dat[3][517][0]=96'h1017a7ee;
sos_loop[0].somModel.sram_ptr[3][517]=3;
sos_loop[0].somModel.sram_dat[3][518][0]=96'h7f128a80;
sos_loop[0].somModel.sram_ptr[3][518]=3;
sos_loop[0].somModel.sram_dat[3][519][0]=96'h7c5925b4;
sos_loop[0].somModel.sram_ptr[3][519]=3;
sos_loop[0].somModel.sram_dat[3][520][0]=96'h4538f048;
sos_loop[0].somModel.sram_ptr[3][520]=3;
sos_loop[0].somModel.sram_dat[3][521][0]=96'ha93c8da7;
sos_loop[0].somModel.sram_ptr[3][521]=3;
sos_loop[0].somModel.sram_dat[3][522][0]=96'hac4a08d6;
sos_loop[0].somModel.sram_ptr[3][522]=3;
sos_loop[0].somModel.sram_dat[3][523][0]=96'h9a0f4cf3;
sos_loop[0].somModel.sram_ptr[3][523]=3;
sos_loop[0].somModel.sram_dat[3][524][0]=96'hf277f763;
sos_loop[0].somModel.sram_ptr[3][524]=3;
sos_loop[0].somModel.sram_dat[3][525][0]=96'h8582cf49;
sos_loop[0].somModel.sram_ptr[3][525]=3;
sos_loop[0].somModel.sram_dat[3][526][0]=96'h93c3f421;
sos_loop[0].somModel.sram_ptr[3][526]=3;
sos_loop[0].somModel.sram_dat[3][527][0]=96'h918c2423;
sos_loop[0].somModel.sram_ptr[3][527]=3;
sos_loop[0].somModel.sram_dat[3][528][0]=96'h9a777ce4;
sos_loop[0].somModel.sram_ptr[3][528]=3;
sos_loop[0].somModel.sram_dat[3][529][0]=96'h36dfd172;
sos_loop[0].somModel.sram_ptr[3][529]=3;
sos_loop[0].somModel.sram_dat[3][530][0]=96'hd5556de3;
sos_loop[0].somModel.sram_ptr[3][530]=3;
sos_loop[0].somModel.sram_dat[3][531][0]=96'hce40b138;
sos_loop[0].somModel.sram_ptr[3][531]=3;
sos_loop[0].somModel.sram_dat[3][532][0]=96'h4aeecfc5;
sos_loop[0].somModel.sram_ptr[3][532]=3;
sos_loop[0].somModel.sram_dat[3][533][0]=96'h3b5012c;
sos_loop[0].somModel.sram_ptr[3][533]=3;
sos_loop[0].somModel.sram_dat[3][534][0]=96'ha397b379;
sos_loop[0].somModel.sram_ptr[3][534]=3;
sos_loop[0].somModel.sram_dat[3][535][0]=96'hc8efbd35;
sos_loop[0].somModel.sram_ptr[3][535]=3;
sos_loop[0].somModel.sram_dat[3][536][0]=96'h197ecb0c;
sos_loop[0].somModel.sram_ptr[3][536]=3;
sos_loop[0].somModel.sram_dat[3][537][0]=96'h3bb510bf;
sos_loop[0].somModel.sram_ptr[3][537]=3;
sos_loop[0].somModel.sram_dat[3][538][0]=96'hc6f6d63e;
sos_loop[0].somModel.sram_ptr[3][538]=3;
sos_loop[0].somModel.sram_dat[3][539][0]=96'h71d6384;
sos_loop[0].somModel.sram_ptr[3][539]=3;
sos_loop[0].somModel.sram_dat[3][540][0]=96'hc552dd1e;
sos_loop[0].somModel.sram_ptr[3][540]=3;
sos_loop[0].somModel.sram_dat[3][541][0]=96'he643bc17;
sos_loop[0].somModel.sram_ptr[3][541]=3;
sos_loop[0].somModel.sram_dat[3][542][0]=96'h43446e4c;
sos_loop[0].somModel.sram_ptr[3][542]=3;
sos_loop[0].somModel.sram_dat[3][543][0]=96'hbcd07cdb;
sos_loop[0].somModel.sram_ptr[3][543]=3;
sos_loop[0].somModel.sram_dat[3][544][0]=96'h7cf14608;
sos_loop[0].somModel.sram_ptr[3][544]=3;
sos_loop[0].somModel.sram_dat[3][545][0]=96'haff02839;
sos_loop[0].somModel.sram_ptr[3][545]=3;
sos_loop[0].somModel.sram_dat[3][546][0]=96'hb6b7b376;
sos_loop[0].somModel.sram_ptr[3][546]=3;
sos_loop[0].somModel.sram_dat[3][547][0]=96'h511eed1;
sos_loop[0].somModel.sram_ptr[3][547]=3;
sos_loop[0].somModel.sram_dat[3][548][0]=96'h6485e04d;
sos_loop[0].somModel.sram_ptr[3][548]=3;
sos_loop[0].somModel.sram_dat[3][549][0]=96'hfb48439e;
sos_loop[0].somModel.sram_ptr[3][549]=3;
sos_loop[0].somModel.sram_dat[3][550][0]=96'h1fb6623a;
sos_loop[0].somModel.sram_ptr[3][550]=3;
sos_loop[0].somModel.sram_dat[3][551][0]=96'h748d035f;
sos_loop[0].somModel.sram_ptr[3][551]=3;
sos_loop[0].somModel.sram_dat[3][552][0]=96'hf999c215;
sos_loop[0].somModel.sram_ptr[3][552]=3;
sos_loop[0].somModel.sram_dat[3][553][0]=96'h36e773ee;
sos_loop[0].somModel.sram_ptr[3][553]=3;
sos_loop[0].somModel.sram_dat[3][554][0]=96'hccdabd4;
sos_loop[0].somModel.sram_ptr[3][554]=3;
sos_loop[0].somModel.sram_dat[3][555][0]=96'hb9bbdeca;
sos_loop[0].somModel.sram_ptr[3][555]=3;
sos_loop[0].somModel.sram_dat[3][556][0]=96'hed764ab2;
sos_loop[0].somModel.sram_ptr[3][556]=3;
sos_loop[0].somModel.sram_dat[3][557][0]=96'h48bac8d7;
sos_loop[0].somModel.sram_ptr[3][557]=3;
sos_loop[0].somModel.sram_dat[3][558][0]=96'h7c5d1f7c;
sos_loop[0].somModel.sram_ptr[3][558]=3;
sos_loop[0].somModel.sram_dat[3][559][0]=96'hb4ce443a;
sos_loop[0].somModel.sram_ptr[3][559]=3;
sos_loop[0].somModel.sram_dat[3][560][0]=96'h65f523a7;
sos_loop[0].somModel.sram_ptr[3][560]=3;
sos_loop[0].somModel.sram_dat[3][561][0]=96'h7875ba6d;
sos_loop[0].somModel.sram_ptr[3][561]=3;
sos_loop[0].somModel.sram_dat[3][562][0]=96'hc13082b4;
sos_loop[0].somModel.sram_ptr[3][562]=3;
sos_loop[0].somModel.sram_dat[3][563][0]=96'hc606c212;
sos_loop[0].somModel.sram_ptr[3][563]=3;
sos_loop[0].somModel.sram_dat[3][564][0]=96'h1e7bb588;
sos_loop[0].somModel.sram_ptr[3][564]=3;
sos_loop[0].somModel.sram_dat[3][565][0]=96'hc05f13a2;
sos_loop[0].somModel.sram_ptr[3][565]=3;
sos_loop[0].somModel.sram_dat[3][566][0]=96'ha10fdd47;
sos_loop[0].somModel.sram_ptr[3][566]=3;
sos_loop[0].somModel.sram_dat[3][567][0]=96'h2cd17cd7;
sos_loop[0].somModel.sram_ptr[3][567]=3;
sos_loop[0].somModel.sram_dat[3][568][0]=96'h116e1259;
sos_loop[0].somModel.sram_ptr[3][568]=3;
sos_loop[0].somModel.sram_dat[3][569][0]=96'h69fd204c;
sos_loop[0].somModel.sram_ptr[3][569]=3;
sos_loop[0].somModel.sram_dat[3][570][0]=96'h12118ecd;
sos_loop[0].somModel.sram_ptr[3][570]=3;
sos_loop[0].somModel.sram_dat[3][571][0]=96'h44d49085;
sos_loop[0].somModel.sram_ptr[3][571]=3;
sos_loop[0].somModel.sram_dat[3][572][0]=96'hd7748be2;
sos_loop[0].somModel.sram_ptr[3][572]=3;
sos_loop[0].somModel.sram_dat[3][573][0]=96'h62dacdb8;
sos_loop[0].somModel.sram_ptr[3][573]=3;
sos_loop[0].somModel.sram_dat[3][574][0]=96'h5d114a9b;
sos_loop[0].somModel.sram_ptr[3][574]=3;
sos_loop[0].somModel.sram_dat[3][575][0]=96'h616bc248;
sos_loop[0].somModel.sram_ptr[3][575]=3;
sos_loop[0].somModel.sram_dat[3][576][0]=96'hb723c38;
sos_loop[0].somModel.sram_ptr[3][576]=3;
sos_loop[0].somModel.sram_dat[3][577][0]=96'hed1fb3c2;
sos_loop[0].somModel.sram_ptr[3][577]=3;
sos_loop[0].somModel.sram_dat[3][578][0]=96'hf845a6c;
sos_loop[0].somModel.sram_ptr[3][578]=3;
sos_loop[0].somModel.sram_dat[3][579][0]=96'hb66c0f85;
sos_loop[0].somModel.sram_ptr[3][579]=3;
sos_loop[0].somModel.sram_dat[3][580][0]=96'hc7600897;
sos_loop[0].somModel.sram_ptr[3][580]=3;
sos_loop[0].somModel.sram_dat[3][581][0]=96'h56100184;
sos_loop[0].somModel.sram_ptr[3][581]=3;
sos_loop[0].somModel.sram_dat[3][582][0]=96'h6bcfe5d6;
sos_loop[0].somModel.sram_ptr[3][582]=3;
sos_loop[0].somModel.sram_dat[3][583][0]=96'hcc94b9b7;
sos_loop[0].somModel.sram_ptr[3][583]=3;
sos_loop[0].somModel.sram_dat[3][584][0]=96'h29e119ed;
sos_loop[0].somModel.sram_ptr[3][584]=3;
sos_loop[0].somModel.sram_dat[3][585][0]=96'he11bfdf4;
sos_loop[0].somModel.sram_ptr[3][585]=3;
sos_loop[0].somModel.sram_dat[3][586][0]=96'h7acacb1f;
sos_loop[0].somModel.sram_ptr[3][586]=3;
sos_loop[0].somModel.sram_dat[3][587][0]=96'hf4956a20;
sos_loop[0].somModel.sram_ptr[3][587]=3;
sos_loop[0].somModel.sram_dat[3][588][0]=96'hd317a971;
sos_loop[0].somModel.sram_ptr[3][588]=3;
sos_loop[0].somModel.sram_dat[3][589][0]=96'h2f31121;
sos_loop[0].somModel.sram_ptr[3][589]=3;
sos_loop[0].somModel.sram_dat[3][590][0]=96'h3e589763;
sos_loop[0].somModel.sram_ptr[3][590]=3;
sos_loop[0].somModel.sram_dat[3][591][0]=96'h5db4743;
sos_loop[0].somModel.sram_ptr[3][591]=3;
sos_loop[0].somModel.sram_dat[3][592][0]=96'hfc1a80cd;
sos_loop[0].somModel.sram_ptr[3][592]=3;
sos_loop[0].somModel.sram_dat[3][593][0]=96'h651ab564;
sos_loop[0].somModel.sram_ptr[3][593]=3;
sos_loop[0].somModel.sram_dat[3][594][0]=96'h8de93c3;
sos_loop[0].somModel.sram_ptr[3][594]=3;
sos_loop[0].somModel.sram_dat[3][595][0]=96'hff37fd0;
sos_loop[0].somModel.sram_ptr[3][595]=3;
sos_loop[0].somModel.sram_dat[3][596][0]=96'h9b657d14;
sos_loop[0].somModel.sram_ptr[3][596]=3;
sos_loop[0].somModel.sram_dat[3][597][0]=96'h6309ce86;
sos_loop[0].somModel.sram_ptr[3][597]=3;
sos_loop[0].somModel.sram_dat[3][598][0]=96'h73716308;
sos_loop[0].somModel.sram_ptr[3][598]=3;
sos_loop[0].somModel.sram_dat[3][599][0]=96'h32c93ff2;
sos_loop[0].somModel.sram_ptr[3][599]=3;
sos_loop[0].somModel.sram_dat[3][600][0]=96'h7883f6d;
sos_loop[0].somModel.sram_ptr[3][600]=3;
sos_loop[0].somModel.sram_dat[3][601][0]=96'hef182c05;
sos_loop[0].somModel.sram_ptr[3][601]=3;
sos_loop[0].somModel.sram_dat[3][602][0]=96'h5cf3d0b;
sos_loop[0].somModel.sram_ptr[3][602]=3;
sos_loop[0].somModel.sram_dat[3][603][0]=96'hfa76e3ad;
sos_loop[0].somModel.sram_ptr[3][603]=3;
sos_loop[0].somModel.sram_dat[3][604][0]=96'hcbd8e504;
sos_loop[0].somModel.sram_ptr[3][604]=3;
sos_loop[0].somModel.sram_dat[3][605][0]=96'h3318e559;
sos_loop[0].somModel.sram_ptr[3][605]=3;
sos_loop[0].somModel.sram_dat[3][606][0]=96'hd2769959;
sos_loop[0].somModel.sram_ptr[3][606]=3;
sos_loop[0].somModel.sram_dat[3][607][0]=96'h54a4165e;
sos_loop[0].somModel.sram_ptr[3][607]=3;
sos_loop[0].somModel.sram_dat[3][608][0]=96'hd19e9f70;
sos_loop[0].somModel.sram_ptr[3][608]=3;
sos_loop[0].somModel.sram_dat[3][609][0]=96'hed963976;
sos_loop[0].somModel.sram_ptr[3][609]=3;
sos_loop[0].somModel.sram_dat[3][610][0]=96'h8c534147;
sos_loop[0].somModel.sram_ptr[3][610]=3;
sos_loop[0].somModel.sram_dat[3][611][0]=96'hd654bf6f;
sos_loop[0].somModel.sram_ptr[3][611]=3;
sos_loop[0].somModel.sram_dat[3][612][0]=96'he8274dc8;
sos_loop[0].somModel.sram_ptr[3][612]=3;
sos_loop[0].somModel.sram_dat[3][613][0]=96'h153e343f;
sos_loop[0].somModel.sram_ptr[3][613]=3;
sos_loop[0].somModel.sram_dat[3][614][0]=96'h76ba647c;
sos_loop[0].somModel.sram_ptr[3][614]=3;
sos_loop[0].somModel.sram_dat[3][615][0]=96'ha78d55ad;
sos_loop[0].somModel.sram_ptr[3][615]=3;
sos_loop[0].somModel.sram_dat[3][616][0]=96'h85bef76c;
sos_loop[0].somModel.sram_ptr[3][616]=3;
sos_loop[0].somModel.sram_dat[3][617][0]=96'h6b8bdd0e;
sos_loop[0].somModel.sram_ptr[3][617]=3;
sos_loop[0].somModel.sram_dat[3][618][0]=96'h3b772627;
sos_loop[0].somModel.sram_ptr[3][618]=3;
sos_loop[0].somModel.sram_dat[3][619][0]=96'h9af419a9;
sos_loop[0].somModel.sram_ptr[3][619]=3;
sos_loop[0].somModel.sram_dat[3][620][0]=96'h33d61638;
sos_loop[0].somModel.sram_ptr[3][620]=3;
sos_loop[0].somModel.sram_dat[3][621][0]=96'he0ce4665;
sos_loop[0].somModel.sram_ptr[3][621]=3;
sos_loop[0].somModel.sram_dat[3][622][0]=96'h1a783a1f;
sos_loop[0].somModel.sram_ptr[3][622]=3;
sos_loop[0].somModel.sram_dat[3][623][0]=96'hc400047;
sos_loop[0].somModel.sram_ptr[3][623]=3;
sos_loop[0].somModel.sram_dat[3][624][0]=96'hefe82a33;
sos_loop[0].somModel.sram_ptr[3][624]=3;
sos_loop[0].somModel.sram_dat[3][625][0]=96'h8fcd729;
sos_loop[0].somModel.sram_ptr[3][625]=3;
sos_loop[0].somModel.sram_dat[3][626][0]=96'h162a2ada;
sos_loop[0].somModel.sram_ptr[3][626]=3;
sos_loop[0].somModel.sram_dat[3][627][0]=96'ha7680901;
sos_loop[0].somModel.sram_ptr[3][627]=3;
sos_loop[0].somModel.sram_dat[3][628][0]=96'h190f7752;
sos_loop[0].somModel.sram_ptr[3][628]=3;
sos_loop[0].somModel.sram_dat[3][629][0]=96'hb6384ac6;
sos_loop[0].somModel.sram_ptr[3][629]=3;
sos_loop[0].somModel.sram_dat[3][630][0]=96'hbbfe5b83;
sos_loop[0].somModel.sram_ptr[3][630]=3;
sos_loop[0].somModel.sram_dat[3][631][0]=96'hcf156c1b;
sos_loop[0].somModel.sram_ptr[3][631]=3;
sos_loop[0].somModel.sram_dat[3][632][0]=96'hda14e4b9;
sos_loop[0].somModel.sram_ptr[3][632]=3;
sos_loop[0].somModel.sram_dat[3][633][0]=96'hf4016e61;
sos_loop[0].somModel.sram_ptr[3][633]=3;
sos_loop[0].somModel.sram_dat[3][634][0]=96'h42f4085d;
sos_loop[0].somModel.sram_ptr[3][634]=3;
sos_loop[0].somModel.sram_dat[3][635][0]=96'h5ea8c2bd;
sos_loop[0].somModel.sram_ptr[3][635]=3;
sos_loop[0].somModel.sram_dat[3][636][0]=96'h303a3b57;
sos_loop[0].somModel.sram_ptr[3][636]=3;
sos_loop[0].somModel.sram_dat[3][637][0]=96'hb7a150b1;
sos_loop[0].somModel.sram_ptr[3][637]=3;
sos_loop[0].somModel.sram_dat[3][638][0]=96'hfb614d0b;
sos_loop[0].somModel.sram_ptr[3][638]=3;
sos_loop[0].somModel.sram_dat[3][639][0]=96'he53edcc3;
sos_loop[0].somModel.sram_ptr[3][639]=3;
sos_loop[0].somModel.sram_dat[3][640][0]=96'h5b0d54c3;
sos_loop[0].somModel.sram_ptr[3][640]=3;
sos_loop[0].somModel.sram_dat[3][641][0]=96'h605ad057;
sos_loop[0].somModel.sram_ptr[3][641]=3;
sos_loop[0].somModel.sram_dat[3][642][0]=96'h8a72fbfe;
sos_loop[0].somModel.sram_ptr[3][642]=3;
sos_loop[0].somModel.sram_dat[3][643][0]=96'h4301aa33;
sos_loop[0].somModel.sram_ptr[3][643]=3;
sos_loop[0].somModel.sram_dat[3][644][0]=96'ha29d6bce;
sos_loop[0].somModel.sram_ptr[3][644]=3;
sos_loop[0].somModel.sram_dat[3][645][0]=96'hc2c68789;
sos_loop[0].somModel.sram_ptr[3][645]=3;
sos_loop[0].somModel.sram_dat[3][646][0]=96'h7370ec2b;
sos_loop[0].somModel.sram_ptr[3][646]=3;
sos_loop[0].somModel.sram_dat[3][647][0]=96'h6989416b;
sos_loop[0].somModel.sram_ptr[3][647]=3;
sos_loop[0].somModel.sram_dat[3][648][0]=96'h6f12824b;
sos_loop[0].somModel.sram_ptr[3][648]=3;
sos_loop[0].somModel.sram_dat[3][649][0]=96'h21ef3f54;
sos_loop[0].somModel.sram_ptr[3][649]=3;
sos_loop[0].somModel.sram_dat[3][650][0]=96'hb9cd2cd9;
sos_loop[0].somModel.sram_ptr[3][650]=3;
sos_loop[0].somModel.sram_dat[3][651][0]=96'hc0e42d17;
sos_loop[0].somModel.sram_ptr[3][651]=3;
sos_loop[0].somModel.sram_dat[3][652][0]=96'h30752c11;
sos_loop[0].somModel.sram_ptr[3][652]=3;
sos_loop[0].somModel.sram_dat[3][653][0]=96'hf36147de;
sos_loop[0].somModel.sram_ptr[3][653]=3;
sos_loop[0].somModel.sram_dat[3][654][0]=96'hdbc68a37;
sos_loop[0].somModel.sram_ptr[3][654]=3;
sos_loop[0].somModel.sram_dat[3][655][0]=96'h77949c5f;
sos_loop[0].somModel.sram_ptr[3][655]=3;
sos_loop[0].somModel.sram_dat[3][656][0]=96'hd4ced086;
sos_loop[0].somModel.sram_ptr[3][656]=3;
sos_loop[0].somModel.sram_dat[3][657][0]=96'hf8b6e64c;
sos_loop[0].somModel.sram_ptr[3][657]=3;
sos_loop[0].somModel.sram_dat[3][658][0]=96'h44618892;
sos_loop[0].somModel.sram_ptr[3][658]=3;
sos_loop[0].somModel.sram_dat[3][659][0]=96'hbcb45bad;
sos_loop[0].somModel.sram_ptr[3][659]=3;
sos_loop[0].somModel.sram_dat[3][660][0]=96'hda6ce781;
sos_loop[0].somModel.sram_ptr[3][660]=3;
sos_loop[0].somModel.sram_dat[3][661][0]=96'hd3268b7;
sos_loop[0].somModel.sram_ptr[3][661]=3;
sos_loop[0].somModel.sram_dat[3][662][0]=96'hb45e9e05;
sos_loop[0].somModel.sram_ptr[3][662]=3;
sos_loop[0].somModel.sram_dat[3][663][0]=96'hcb3466e1;
sos_loop[0].somModel.sram_ptr[3][663]=3;
sos_loop[0].somModel.sram_dat[3][664][0]=96'h343705e1;
sos_loop[0].somModel.sram_ptr[3][664]=3;
sos_loop[0].somModel.sram_dat[3][665][0]=96'hf235af9a;
sos_loop[0].somModel.sram_ptr[3][665]=3;
sos_loop[0].somModel.sram_dat[3][666][0]=96'h740ad0a0;
sos_loop[0].somModel.sram_ptr[3][666]=3;
sos_loop[0].somModel.sram_dat[3][667][0]=96'he7680fcb;
sos_loop[0].somModel.sram_ptr[3][667]=3;
sos_loop[0].somModel.sram_dat[3][668][0]=96'hd1ea0b9b;
sos_loop[0].somModel.sram_ptr[3][668]=3;
sos_loop[0].somModel.sram_dat[3][669][0]=96'h4e15f57c;
sos_loop[0].somModel.sram_ptr[3][669]=3;
sos_loop[0].somModel.sram_dat[3][670][0]=96'hc059765f;
sos_loop[0].somModel.sram_ptr[3][670]=3;
sos_loop[0].somModel.sram_dat[3][671][0]=96'h9df097da;
sos_loop[0].somModel.sram_ptr[3][671]=3;
sos_loop[0].somModel.sram_dat[3][672][0]=96'hc6549881;
sos_loop[0].somModel.sram_ptr[3][672]=3;
sos_loop[0].somModel.sram_dat[3][673][0]=96'h895b90ac;
sos_loop[0].somModel.sram_ptr[3][673]=3;
sos_loop[0].somModel.sram_dat[3][674][0]=96'h41466398;
sos_loop[0].somModel.sram_ptr[3][674]=3;
sos_loop[0].somModel.sram_dat[3][675][0]=96'hc6a8e81e;
sos_loop[0].somModel.sram_ptr[3][675]=3;
sos_loop[0].somModel.sram_dat[3][676][0]=96'h93ab9460;
sos_loop[0].somModel.sram_ptr[3][676]=3;
sos_loop[0].somModel.sram_dat[3][677][0]=96'he90e7140;
sos_loop[0].somModel.sram_ptr[3][677]=3;
sos_loop[0].somModel.sram_dat[3][678][0]=96'hf8fb4acb;
sos_loop[0].somModel.sram_ptr[3][678]=3;
sos_loop[0].somModel.sram_dat[3][679][0]=96'h1031b5dd;
sos_loop[0].somModel.sram_ptr[3][679]=3;
sos_loop[0].somModel.sram_dat[3][680][0]=96'he4dc251b;
sos_loop[0].somModel.sram_ptr[3][680]=3;
sos_loop[0].somModel.sram_dat[3][681][0]=96'h53d482fa;
sos_loop[0].somModel.sram_ptr[3][681]=3;
sos_loop[0].somModel.sram_dat[3][682][0]=96'he0ff78f3;
sos_loop[0].somModel.sram_ptr[3][682]=3;
sos_loop[0].somModel.sram_dat[3][683][0]=96'h1af2f077;
sos_loop[0].somModel.sram_ptr[3][683]=3;
sos_loop[0].somModel.sram_dat[3][684][0]=96'h7bdb5913;
sos_loop[0].somModel.sram_ptr[3][684]=3;
sos_loop[0].somModel.sram_dat[3][685][0]=96'h8f40dddc;
sos_loop[0].somModel.sram_ptr[3][685]=3;
sos_loop[0].somModel.sram_dat[3][686][0]=96'h17f3c692;
sos_loop[0].somModel.sram_ptr[3][686]=3;
sos_loop[0].somModel.sram_dat[3][687][0]=96'h75db959a;
sos_loop[0].somModel.sram_ptr[3][687]=3;
sos_loop[0].somModel.sram_dat[3][688][0]=96'h755727cf;
sos_loop[0].somModel.sram_ptr[3][688]=3;
sos_loop[0].somModel.sram_dat[3][689][0]=96'h374bbaf3;
sos_loop[0].somModel.sram_ptr[3][689]=3;
sos_loop[0].somModel.sram_dat[3][690][0]=96'h8a7eca48;
sos_loop[0].somModel.sram_ptr[3][690]=3;
sos_loop[0].somModel.sram_dat[3][691][0]=96'h75d671e7;
sos_loop[0].somModel.sram_ptr[3][691]=3;
sos_loop[0].somModel.sram_dat[3][692][0]=96'hf026b004;
sos_loop[0].somModel.sram_ptr[3][692]=3;
sos_loop[0].somModel.sram_dat[3][693][0]=96'hd482915d;
sos_loop[0].somModel.sram_ptr[3][693]=3;
sos_loop[0].somModel.sram_dat[3][694][0]=96'hee8ec632;
sos_loop[0].somModel.sram_ptr[3][694]=3;
sos_loop[0].somModel.sram_dat[3][695][0]=96'h2a2556b1;
sos_loop[0].somModel.sram_ptr[3][695]=3;
sos_loop[0].somModel.sram_dat[3][696][0]=96'h3aa3da2c;
sos_loop[0].somModel.sram_ptr[3][696]=3;
sos_loop[0].somModel.sram_dat[3][697][0]=96'h62e599fd;
sos_loop[0].somModel.sram_ptr[3][697]=3;
sos_loop[0].somModel.sram_dat[3][698][0]=96'h3ad006a9;
sos_loop[0].somModel.sram_ptr[3][698]=3;
sos_loop[0].somModel.sram_dat[3][699][0]=96'hf129a13;
sos_loop[0].somModel.sram_ptr[3][699]=3;
sos_loop[0].somModel.sram_dat[3][700][0]=96'hbd3eb75c;
sos_loop[0].somModel.sram_ptr[3][700]=3;
sos_loop[0].somModel.cfg_tbl_sel[3] = 3;
sos_loop[0].somModel.cfg_dat_sel[3] = 1;
sos_loop[0].somModel.cfg_dat_vld[3] = 1;
sos_loop[0].somModel.cfg_miss_ptr[3] = 0;
sos_loop[0].somModel.tcam_data[4][0][0]=80'h00000000000000000000;
sos_loop[0].somModel.tcam_mask[4][0][0]=80'hffffffffffffffffffff;
sos_loop[0].somModel.tcam_data[4][1][0]=80'h000000000000007f1ea9;
sos_loop[0].somModel.tcam_mask[4][1][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][2][0]=80'h0000000000000018d7d4;
sos_loop[0].somModel.tcam_mask[4][2][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][3][0]=80'h00000000000000879503;
sos_loop[0].somModel.tcam_mask[4][3][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][4][0]=80'h00000000000000795e9d;
sos_loop[0].somModel.tcam_mask[4][4][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][5][0]=80'h00000000000000d8811f;
sos_loop[0].somModel.tcam_mask[4][5][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][6][0]=80'h00000000000000f72c4f;
sos_loop[0].somModel.tcam_mask[4][6][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][7][0]=80'h0000000000000045bc37;
sos_loop[0].somModel.tcam_mask[4][7][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][8][0]=80'h00000000000000a9ca1e;
sos_loop[0].somModel.tcam_mask[4][8][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][9][0]=80'h0000000000000095fadc;
sos_loop[0].somModel.tcam_mask[4][9][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][10][0]=80'h00000000000000fd7856;
sos_loop[0].somModel.tcam_mask[4][10][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][11][0]=80'h000000000000003ac1d0;
sos_loop[0].somModel.tcam_mask[4][11][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][12][0]=80'h000000000000000c47e0;
sos_loop[0].somModel.tcam_mask[4][12][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][13][0]=80'h00000000000000fb27f9;
sos_loop[0].somModel.tcam_mask[4][13][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][14][0]=80'h0000000000000018fca4;
sos_loop[0].somModel.tcam_mask[4][14][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][15][0]=80'h000000000000002e4356;
sos_loop[0].somModel.tcam_mask[4][15][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][16][0]=80'h0000000000000056a40c;
sos_loop[0].somModel.tcam_mask[4][16][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][17][0]=80'h0000000000000018540e;
sos_loop[0].somModel.tcam_mask[4][17][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][18][0]=80'h00000000000000ea2b44;
sos_loop[0].somModel.tcam_mask[4][18][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][19][0]=80'h0000000000000084c769;
sos_loop[0].somModel.tcam_mask[4][19][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][20][0]=80'h000000000000009ae0b9;
sos_loop[0].somModel.tcam_mask[4][20][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][21][0]=80'h00000000000000a15356;
sos_loop[0].somModel.tcam_mask[4][21][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][22][0]=80'h000000000000005a0605;
sos_loop[0].somModel.tcam_mask[4][22][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][23][0]=80'h000000000000006fe0cb;
sos_loop[0].somModel.tcam_mask[4][23][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][24][0]=80'h00000000000000e646d6;
sos_loop[0].somModel.tcam_mask[4][24][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][25][0]=80'h000000000000000a2d6b;
sos_loop[0].somModel.tcam_mask[4][25][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][26][0]=80'h00000000000000f04d5b;
sos_loop[0].somModel.tcam_mask[4][26][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][27][0]=80'h000000000000004c578c;
sos_loop[0].somModel.tcam_mask[4][27][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][28][0]=80'h00000000000000888d1f;
sos_loop[0].somModel.tcam_mask[4][28][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][29][0]=80'h000000000000002ca3fe;
sos_loop[0].somModel.tcam_mask[4][29][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][30][0]=80'h0000000000000063455b;
sos_loop[0].somModel.tcam_mask[4][30][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][31][0]=80'h000000000000002768c3;
sos_loop[0].somModel.tcam_mask[4][31][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][32][0]=80'h000000000000007cb8cb;
sos_loop[0].somModel.tcam_mask[4][32][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][33][0]=80'h0000000000000062f735;
sos_loop[0].somModel.tcam_mask[4][33][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][34][0]=80'h000000000000002fa2ac;
sos_loop[0].somModel.tcam_mask[4][34][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][35][0]=80'h000000000000006b0b30;
sos_loop[0].somModel.tcam_mask[4][35][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][36][0]=80'h00000000000000dc4120;
sos_loop[0].somModel.tcam_mask[4][36][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][37][0]=80'h00000000000000d471aa;
sos_loop[0].somModel.tcam_mask[4][37][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][38][0]=80'h0000000000000040a7fc;
sos_loop[0].somModel.tcam_mask[4][38][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][39][0]=80'h00000000000000ac33c6;
sos_loop[0].somModel.tcam_mask[4][39][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][40][0]=80'h00000000000000109775;
sos_loop[0].somModel.tcam_mask[4][40][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][41][0]=80'h00000000000000c3ff40;
sos_loop[0].somModel.tcam_mask[4][41][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][42][0]=80'h00000000000000283e24;
sos_loop[0].somModel.tcam_mask[4][42][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][43][0]=80'h00000000000000d2bca2;
sos_loop[0].somModel.tcam_mask[4][43][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][44][0]=80'h000000000000005178a5;
sos_loop[0].somModel.tcam_mask[4][44][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][45][0]=80'h000000000000009ab1a5;
sos_loop[0].somModel.tcam_mask[4][45][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][46][0]=80'h00000000000000dd0418;
sos_loop[0].somModel.tcam_mask[4][46][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][47][0]=80'h000000000000004341e8;
sos_loop[0].somModel.tcam_mask[4][47][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][48][0]=80'h00000000000000beafd2;
sos_loop[0].somModel.tcam_mask[4][48][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][49][0]=80'h00000000000000653c68;
sos_loop[0].somModel.tcam_mask[4][49][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][50][0]=80'h00000000000000c2f7fb;
sos_loop[0].somModel.tcam_mask[4][50][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][51][0]=80'h000000000000002ec425;
sos_loop[0].somModel.tcam_mask[4][51][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][52][0]=80'h0000000000000039f1b8;
sos_loop[0].somModel.tcam_mask[4][52][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][53][0]=80'h0000000000000065b81f;
sos_loop[0].somModel.tcam_mask[4][53][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][54][0]=80'h00000000000000e84bff;
sos_loop[0].somModel.tcam_mask[4][54][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][55][0]=80'h000000000000006f12c1;
sos_loop[0].somModel.tcam_mask[4][55][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][56][0]=80'h00000000000000638539;
sos_loop[0].somModel.tcam_mask[4][56][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][57][0]=80'h0000000000000074386b;
sos_loop[0].somModel.tcam_mask[4][57][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][58][0]=80'h000000000000006ec296;
sos_loop[0].somModel.tcam_mask[4][58][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][59][0]=80'h000000000000009dc45a;
sos_loop[0].somModel.tcam_mask[4][59][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][60][0]=80'h000000000000007bdeb2;
sos_loop[0].somModel.tcam_mask[4][60][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][61][0]=80'h00000000000000109400;
sos_loop[0].somModel.tcam_mask[4][61][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][62][0]=80'h000000000000003ed34b;
sos_loop[0].somModel.tcam_mask[4][62][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][63][0]=80'h0000000000000083a39a;
sos_loop[0].somModel.tcam_mask[4][63][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][64][0]=80'h00000000000000b39350;
sos_loop[0].somModel.tcam_mask[4][64][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][65][0]=80'h000000000000003fd68e;
sos_loop[0].somModel.tcam_mask[4][65][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][66][0]=80'h00000000000000168dc8;
sos_loop[0].somModel.tcam_mask[4][66][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][67][0]=80'h00000000000000c7d864;
sos_loop[0].somModel.tcam_mask[4][67][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][68][0]=80'h000000000000006ac4b8;
sos_loop[0].somModel.tcam_mask[4][68][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][69][0]=80'h0000000000000029c5fa;
sos_loop[0].somModel.tcam_mask[4][69][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][70][0]=80'h000000000000007775e4;
sos_loop[0].somModel.tcam_mask[4][70][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][71][0]=80'h00000000000000354a38;
sos_loop[0].somModel.tcam_mask[4][71][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][72][0]=80'h00000000000000482f82;
sos_loop[0].somModel.tcam_mask[4][72][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][73][0]=80'h000000000000008f4dc7;
sos_loop[0].somModel.tcam_mask[4][73][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][74][0]=80'h000000000000002f794e;
sos_loop[0].somModel.tcam_mask[4][74][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][75][0]=80'h00000000000000c688bd;
sos_loop[0].somModel.tcam_mask[4][75][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][76][0]=80'h000000000000008c6bf8;
sos_loop[0].somModel.tcam_mask[4][76][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][77][0]=80'h000000000000004a580d;
sos_loop[0].somModel.tcam_mask[4][77][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][78][0]=80'h00000000000000e51d07;
sos_loop[0].somModel.tcam_mask[4][78][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][79][0]=80'h000000000000006576cb;
sos_loop[0].somModel.tcam_mask[4][79][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][80][0]=80'h00000000000000672b33;
sos_loop[0].somModel.tcam_mask[4][80][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][81][0]=80'h00000000000000765369;
sos_loop[0].somModel.tcam_mask[4][81][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][82][0]=80'h00000000000000065548;
sos_loop[0].somModel.tcam_mask[4][82][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][83][0]=80'h00000000000000fa8b7f;
sos_loop[0].somModel.tcam_mask[4][83][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][84][0]=80'h000000000000009e0149;
sos_loop[0].somModel.tcam_mask[4][84][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][85][0]=80'h000000000000003700bc;
sos_loop[0].somModel.tcam_mask[4][85][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][86][0]=80'h00000000000000a26d54;
sos_loop[0].somModel.tcam_mask[4][86][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][87][0]=80'h00000000000000485e50;
sos_loop[0].somModel.tcam_mask[4][87][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][88][0]=80'h000000000000004e377c;
sos_loop[0].somModel.tcam_mask[4][88][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][89][0]=80'h00000000000000290bd8;
sos_loop[0].somModel.tcam_mask[4][89][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][90][0]=80'h0000000000000079eac3;
sos_loop[0].somModel.tcam_mask[4][90][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][91][0]=80'h00000000000000aeb963;
sos_loop[0].somModel.tcam_mask[4][91][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][92][0]=80'h000000000000000e60f6;
sos_loop[0].somModel.tcam_mask[4][92][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][93][0]=80'h00000000000000ebc64c;
sos_loop[0].somModel.tcam_mask[4][93][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][94][0]=80'h00000000000000fd79da;
sos_loop[0].somModel.tcam_mask[4][94][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][95][0]=80'h000000000000005f903f;
sos_loop[0].somModel.tcam_mask[4][95][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][96][0]=80'h000000000000008c6098;
sos_loop[0].somModel.tcam_mask[4][96][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][97][0]=80'h0000000000000052bbf8;
sos_loop[0].somModel.tcam_mask[4][97][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][98][0]=80'h0000000000000067064a;
sos_loop[0].somModel.tcam_mask[4][98][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][99][0]=80'h00000000000000eda0ac;
sos_loop[0].somModel.tcam_mask[4][99][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][100][0]=80'h000000000000009fe0b2;
sos_loop[0].somModel.tcam_mask[4][100][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][101][0]=80'h000000000000002b0b9e;
sos_loop[0].somModel.tcam_mask[4][101][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][102][0]=80'h000000000000008ed315;
sos_loop[0].somModel.tcam_mask[4][102][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][103][0]=80'h000000000000003fa5eb;
sos_loop[0].somModel.tcam_mask[4][103][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][104][0]=80'h00000000000000d5a9ea;
sos_loop[0].somModel.tcam_mask[4][104][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][105][0]=80'h000000000000003b5063;
sos_loop[0].somModel.tcam_mask[4][105][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][106][0]=80'h000000000000003de498;
sos_loop[0].somModel.tcam_mask[4][106][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][107][0]=80'h0000000000000034d05b;
sos_loop[0].somModel.tcam_mask[4][107][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][108][0]=80'h000000000000009906b4;
sos_loop[0].somModel.tcam_mask[4][108][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][109][0]=80'h000000000000008e8559;
sos_loop[0].somModel.tcam_mask[4][109][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][110][0]=80'h000000000000000e3f52;
sos_loop[0].somModel.tcam_mask[4][110][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][111][0]=80'h000000000000004b4571;
sos_loop[0].somModel.tcam_mask[4][111][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][112][0]=80'h000000000000001da95e;
sos_loop[0].somModel.tcam_mask[4][112][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][113][0]=80'h00000000000000f8a77d;
sos_loop[0].somModel.tcam_mask[4][113][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][114][0]=80'h000000000000000773e7;
sos_loop[0].somModel.tcam_mask[4][114][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][115][0]=80'h00000000000000cc18d8;
sos_loop[0].somModel.tcam_mask[4][115][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][116][0]=80'h00000000000000523f2c;
sos_loop[0].somModel.tcam_mask[4][116][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][117][0]=80'h00000000000000d32eb1;
sos_loop[0].somModel.tcam_mask[4][117][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][118][0]=80'h00000000000000b10a04;
sos_loop[0].somModel.tcam_mask[4][118][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][119][0]=80'h000000000000009e289a;
sos_loop[0].somModel.tcam_mask[4][119][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][120][0]=80'h000000000000003f745c;
sos_loop[0].somModel.tcam_mask[4][120][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][121][0]=80'h00000000000000b4d716;
sos_loop[0].somModel.tcam_mask[4][121][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][122][0]=80'h00000000000000353aba;
sos_loop[0].somModel.tcam_mask[4][122][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][123][0]=80'h00000000000000138266;
sos_loop[0].somModel.tcam_mask[4][123][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][124][0]=80'h0000000000000098c3a8;
sos_loop[0].somModel.tcam_mask[4][124][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][125][0]=80'h00000000000000a72bb0;
sos_loop[0].somModel.tcam_mask[4][125][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][126][0]=80'h00000000000000f0a808;
sos_loop[0].somModel.tcam_mask[4][126][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][127][0]=80'h000000000000002ecc7c;
sos_loop[0].somModel.tcam_mask[4][127][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][128][0]=80'h0000000000000070432e;
sos_loop[0].somModel.tcam_mask[4][128][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][129][0]=80'h000000000000009e5629;
sos_loop[0].somModel.tcam_mask[4][129][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][130][0]=80'h00000000000000b9028f;
sos_loop[0].somModel.tcam_mask[4][130][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][131][0]=80'h000000000000007d192f;
sos_loop[0].somModel.tcam_mask[4][131][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][132][0]=80'h000000000000009f9291;
sos_loop[0].somModel.tcam_mask[4][132][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][133][0]=80'h00000000000000ee6a20;
sos_loop[0].somModel.tcam_mask[4][133][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][134][0]=80'h0000000000000053672d;
sos_loop[0].somModel.tcam_mask[4][134][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][135][0]=80'h00000000000000dd027c;
sos_loop[0].somModel.tcam_mask[4][135][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][136][0]=80'h000000000000000dc08c;
sos_loop[0].somModel.tcam_mask[4][136][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][137][0]=80'h0000000000000058402c;
sos_loop[0].somModel.tcam_mask[4][137][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][138][0]=80'h00000000000000c81a4a;
sos_loop[0].somModel.tcam_mask[4][138][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][139][0]=80'h00000000000000edd5d3;
sos_loop[0].somModel.tcam_mask[4][139][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][140][0]=80'h00000000000000004b52;
sos_loop[0].somModel.tcam_mask[4][140][0]=80'hffffffffffffffff8000;
sos_loop[0].somModel.tcam_data[4][141][0]=80'h00000000000000e03ed4;
sos_loop[0].somModel.tcam_mask[4][141][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][142][0]=80'h000000000000007e9436;
sos_loop[0].somModel.tcam_mask[4][142][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][143][0]=80'h00000000000000784bef;
sos_loop[0].somModel.tcam_mask[4][143][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][144][0]=80'h0000000000000042f39d;
sos_loop[0].somModel.tcam_mask[4][144][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][145][0]=80'h00000000000000be6a7e;
sos_loop[0].somModel.tcam_mask[4][145][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][146][0]=80'h00000000000000826f57;
sos_loop[0].somModel.tcam_mask[4][146][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][147][0]=80'h00000000000000029e2c;
sos_loop[0].somModel.tcam_mask[4][147][0]=80'hfffffffffffffffc0000;
sos_loop[0].somModel.tcam_data[4][148][0]=80'h0000000000000029c960;
sos_loop[0].somModel.tcam_mask[4][148][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][149][0]=80'h0000000000000019c756;
sos_loop[0].somModel.tcam_mask[4][149][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][150][0]=80'h0000000000000001fbdf;
sos_loop[0].somModel.tcam_mask[4][150][0]=80'hfffffffffffffffe0000;
sos_loop[0].somModel.tcam_data[4][151][0]=80'h000000000000000798a3;
sos_loop[0].somModel.tcam_mask[4][151][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][152][0]=80'h00000000000000376c99;
sos_loop[0].somModel.tcam_mask[4][152][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][153][0]=80'h000000000000002e7c93;
sos_loop[0].somModel.tcam_mask[4][153][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][154][0]=80'h000000000000006e0c48;
sos_loop[0].somModel.tcam_mask[4][154][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][155][0]=80'h000000000000007848e4;
sos_loop[0].somModel.tcam_mask[4][155][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][156][0]=80'h00000000000000eab49b;
sos_loop[0].somModel.tcam_mask[4][156][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][157][0]=80'h000000000000003c4183;
sos_loop[0].somModel.tcam_mask[4][157][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][158][0]=80'h00000000000000206e77;
sos_loop[0].somModel.tcam_mask[4][158][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][159][0]=80'h0000000000000060af7b;
sos_loop[0].somModel.tcam_mask[4][159][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][160][0]=80'h00000000000000532847;
sos_loop[0].somModel.tcam_mask[4][160][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][161][0]=80'h00000000000000bad608;
sos_loop[0].somModel.tcam_mask[4][161][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][162][0]=80'h0000000000000047a19a;
sos_loop[0].somModel.tcam_mask[4][162][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][163][0]=80'h00000000000000f8c422;
sos_loop[0].somModel.tcam_mask[4][163][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][164][0]=80'h000000000000009c50ab;
sos_loop[0].somModel.tcam_mask[4][164][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][165][0]=80'h000000000000002c4a16;
sos_loop[0].somModel.tcam_mask[4][165][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][166][0]=80'h00000000000000e2f212;
sos_loop[0].somModel.tcam_mask[4][166][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][167][0]=80'h0000000000000032b6e2;
sos_loop[0].somModel.tcam_mask[4][167][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][168][0]=80'h00000000000000501cd9;
sos_loop[0].somModel.tcam_mask[4][168][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][169][0]=80'h0000000000000059d817;
sos_loop[0].somModel.tcam_mask[4][169][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][170][0]=80'h0000000000000079c4b3;
sos_loop[0].somModel.tcam_mask[4][170][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][171][0]=80'h00000000000000dbfb38;
sos_loop[0].somModel.tcam_mask[4][171][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][172][0]=80'h000000000000003c8d91;
sos_loop[0].somModel.tcam_mask[4][172][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][173][0]=80'h00000000000000700b97;
sos_loop[0].somModel.tcam_mask[4][173][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][174][0]=80'h000000000000006a6798;
sos_loop[0].somModel.tcam_mask[4][174][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][175][0]=80'h00000000000000b16541;
sos_loop[0].somModel.tcam_mask[4][175][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][176][0]=80'h00000000000000148fdc;
sos_loop[0].somModel.tcam_mask[4][176][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][177][0]=80'h00000000000000c77ae0;
sos_loop[0].somModel.tcam_mask[4][177][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][178][0]=80'h00000000000000289a41;
sos_loop[0].somModel.tcam_mask[4][178][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][179][0]=80'h00000000000000cce9c6;
sos_loop[0].somModel.tcam_mask[4][179][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][180][0]=80'h000000000000003293d0;
sos_loop[0].somModel.tcam_mask[4][180][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][181][0]=80'h0000000000000085fe27;
sos_loop[0].somModel.tcam_mask[4][181][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][182][0]=80'h000000000000007de321;
sos_loop[0].somModel.tcam_mask[4][182][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][183][0]=80'h00000000000000556878;
sos_loop[0].somModel.tcam_mask[4][183][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][184][0]=80'h00000000000000a2e200;
sos_loop[0].somModel.tcam_mask[4][184][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][185][0]=80'h00000000000000f7b199;
sos_loop[0].somModel.tcam_mask[4][185][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][186][0]=80'h000000000000004e7d0f;
sos_loop[0].somModel.tcam_mask[4][186][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][187][0]=80'h000000000000002932d5;
sos_loop[0].somModel.tcam_mask[4][187][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][188][0]=80'h00000000000000f10ee2;
sos_loop[0].somModel.tcam_mask[4][188][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][189][0]=80'h00000000000000d3cb30;
sos_loop[0].somModel.tcam_mask[4][189][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][190][0]=80'h00000000000000dc4082;
sos_loop[0].somModel.tcam_mask[4][190][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][191][0]=80'h000000000000004680df;
sos_loop[0].somModel.tcam_mask[4][191][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][192][0]=80'h000000000000003e3ace;
sos_loop[0].somModel.tcam_mask[4][192][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][193][0]=80'h00000000000000278237;
sos_loop[0].somModel.tcam_mask[4][193][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][194][0]=80'h00000000000000f58b4b;
sos_loop[0].somModel.tcam_mask[4][194][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][195][0]=80'h0000000000000053a60b;
sos_loop[0].somModel.tcam_mask[4][195][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][196][0]=80'h0000000000000029bce4;
sos_loop[0].somModel.tcam_mask[4][196][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][197][0]=80'h00000000000000bf1a0a;
sos_loop[0].somModel.tcam_mask[4][197][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][198][0]=80'h00000000000000e19318;
sos_loop[0].somModel.tcam_mask[4][198][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][199][0]=80'h0000000000000044d266;
sos_loop[0].somModel.tcam_mask[4][199][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][200][0]=80'h00000000000000a6b455;
sos_loop[0].somModel.tcam_mask[4][200][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][201][0]=80'h00000000000000a1ed9d;
sos_loop[0].somModel.tcam_mask[4][201][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][202][0]=80'h000000000000004fc0f7;
sos_loop[0].somModel.tcam_mask[4][202][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][203][0]=80'h0000000000000083eaaf;
sos_loop[0].somModel.tcam_mask[4][203][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][204][0]=80'h0000000000000001d8f2;
sos_loop[0].somModel.tcam_mask[4][204][0]=80'hfffffffffffffffe0000;
sos_loop[0].somModel.tcam_data[4][205][0]=80'h000000000000000c8461;
sos_loop[0].somModel.tcam_mask[4][205][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][206][0]=80'h000000000000005a9ad8;
sos_loop[0].somModel.tcam_mask[4][206][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][207][0]=80'h0000000000000045adc4;
sos_loop[0].somModel.tcam_mask[4][207][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][208][0]=80'h0000000000000044e7f5;
sos_loop[0].somModel.tcam_mask[4][208][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][209][0]=80'h000000000000004a5dba;
sos_loop[0].somModel.tcam_mask[4][209][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][210][0]=80'h0000000000000082d37a;
sos_loop[0].somModel.tcam_mask[4][210][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][211][0]=80'h00000000000000a5936e;
sos_loop[0].somModel.tcam_mask[4][211][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][212][0]=80'h0000000000000007b239;
sos_loop[0].somModel.tcam_mask[4][212][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][213][0]=80'h0000000000000012fd45;
sos_loop[0].somModel.tcam_mask[4][213][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][214][0]=80'h00000000000000842ec1;
sos_loop[0].somModel.tcam_mask[4][214][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][215][0]=80'h000000000000005fee07;
sos_loop[0].somModel.tcam_mask[4][215][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][216][0]=80'h00000000000000386dc0;
sos_loop[0].somModel.tcam_mask[4][216][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][217][0]=80'h0000000000000030a003;
sos_loop[0].somModel.tcam_mask[4][217][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][218][0]=80'h0000000000000069dabf;
sos_loop[0].somModel.tcam_mask[4][218][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][219][0]=80'h000000000000000c8cd9;
sos_loop[0].somModel.tcam_mask[4][219][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][220][0]=80'h0000000000000020926d;
sos_loop[0].somModel.tcam_mask[4][220][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][221][0]=80'h00000000000000c358af;
sos_loop[0].somModel.tcam_mask[4][221][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][222][0]=80'h000000000000005bb9eb;
sos_loop[0].somModel.tcam_mask[4][222][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][223][0]=80'h00000000000000b1e73e;
sos_loop[0].somModel.tcam_mask[4][223][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][224][0]=80'h00000000000000591f46;
sos_loop[0].somModel.tcam_mask[4][224][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][225][0]=80'h000000000000007367d3;
sos_loop[0].somModel.tcam_mask[4][225][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][226][0]=80'h00000000000000638b62;
sos_loop[0].somModel.tcam_mask[4][226][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][227][0]=80'h00000000000000637b90;
sos_loop[0].somModel.tcam_mask[4][227][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][228][0]=80'h000000000000008d74b6;
sos_loop[0].somModel.tcam_mask[4][228][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][229][0]=80'h000000000000005c8f52;
sos_loop[0].somModel.tcam_mask[4][229][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][230][0]=80'h00000000000000d7ee49;
sos_loop[0].somModel.tcam_mask[4][230][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][231][0]=80'h00000000000000d72b91;
sos_loop[0].somModel.tcam_mask[4][231][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][232][0]=80'h00000000000000816c24;
sos_loop[0].somModel.tcam_mask[4][232][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][233][0]=80'h00000000000000de97a8;
sos_loop[0].somModel.tcam_mask[4][233][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][234][0]=80'h000000000000004ef26b;
sos_loop[0].somModel.tcam_mask[4][234][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][235][0]=80'h00000000000000afbc7c;
sos_loop[0].somModel.tcam_mask[4][235][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][236][0]=80'h00000000000000337d7d;
sos_loop[0].somModel.tcam_mask[4][236][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][237][0]=80'h00000000000000781a2b;
sos_loop[0].somModel.tcam_mask[4][237][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][238][0]=80'h00000000000000b4e99c;
sos_loop[0].somModel.tcam_mask[4][238][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][239][0]=80'h00000000000000a1d931;
sos_loop[0].somModel.tcam_mask[4][239][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][240][0]=80'h000000000000002e3027;
sos_loop[0].somModel.tcam_mask[4][240][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][241][0]=80'h00000000000000f983f9;
sos_loop[0].somModel.tcam_mask[4][241][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][242][0]=80'h0000000000000056ed80;
sos_loop[0].somModel.tcam_mask[4][242][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][243][0]=80'h000000000000005200ab;
sos_loop[0].somModel.tcam_mask[4][243][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][244][0]=80'h00000000000000637797;
sos_loop[0].somModel.tcam_mask[4][244][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][245][0]=80'h00000000000000dd2137;
sos_loop[0].somModel.tcam_mask[4][245][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][246][0]=80'h00000000000000fd2416;
sos_loop[0].somModel.tcam_mask[4][246][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][247][0]=80'h00000000000000f3a4f0;
sos_loop[0].somModel.tcam_mask[4][247][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][248][0]=80'h0000000000000044c886;
sos_loop[0].somModel.tcam_mask[4][248][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][249][0]=80'h00000000000000ceb410;
sos_loop[0].somModel.tcam_mask[4][249][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][250][0]=80'h00000000000000f59b12;
sos_loop[0].somModel.tcam_mask[4][250][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][251][0]=80'h00000000000000e49bd0;
sos_loop[0].somModel.tcam_mask[4][251][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][252][0]=80'h00000000000000638997;
sos_loop[0].somModel.tcam_mask[4][252][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][253][0]=80'h000000000000002f7580;
sos_loop[0].somModel.tcam_mask[4][253][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][254][0]=80'h000000000000001c10a8;
sos_loop[0].somModel.tcam_mask[4][254][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][255][0]=80'h00000000000000879f04;
sos_loop[0].somModel.tcam_mask[4][255][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][256][0]=80'h00000000000000bab2c4;
sos_loop[0].somModel.tcam_mask[4][256][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][257][0]=80'h00000000000000a22715;
sos_loop[0].somModel.tcam_mask[4][257][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][258][0]=80'h00000000000000f23b5e;
sos_loop[0].somModel.tcam_mask[4][258][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][259][0]=80'h00000000000000fdc001;
sos_loop[0].somModel.tcam_mask[4][259][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][260][0]=80'h00000000000000288bf0;
sos_loop[0].somModel.tcam_mask[4][260][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][261][0]=80'h00000000000000662d40;
sos_loop[0].somModel.tcam_mask[4][261][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][262][0]=80'h0000000000000072cef9;
sos_loop[0].somModel.tcam_mask[4][262][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][263][0]=80'h00000000000000087666;
sos_loop[0].somModel.tcam_mask[4][263][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][264][0]=80'h00000000000000f522c4;
sos_loop[0].somModel.tcam_mask[4][264][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][265][0]=80'h00000000000000cf63c5;
sos_loop[0].somModel.tcam_mask[4][265][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][266][0]=80'h00000000000000e18e89;
sos_loop[0].somModel.tcam_mask[4][266][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][267][0]=80'h00000000000000a2bc46;
sos_loop[0].somModel.tcam_mask[4][267][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][268][0]=80'h0000000000000041996f;
sos_loop[0].somModel.tcam_mask[4][268][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][269][0]=80'h000000000000005e2a51;
sos_loop[0].somModel.tcam_mask[4][269][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][270][0]=80'h0000000000000046b451;
sos_loop[0].somModel.tcam_mask[4][270][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][271][0]=80'h00000000000000ee2aae;
sos_loop[0].somModel.tcam_mask[4][271][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][272][0]=80'h00000000000000b33948;
sos_loop[0].somModel.tcam_mask[4][272][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][273][0]=80'h000000000000007587fe;
sos_loop[0].somModel.tcam_mask[4][273][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][274][0]=80'h000000000000004584c5;
sos_loop[0].somModel.tcam_mask[4][274][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][275][0]=80'h000000000000004532c5;
sos_loop[0].somModel.tcam_mask[4][275][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][276][0]=80'h000000000000007754d8;
sos_loop[0].somModel.tcam_mask[4][276][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][277][0]=80'h0000000000000002b77b;
sos_loop[0].somModel.tcam_mask[4][277][0]=80'hfffffffffffffffc0000;
sos_loop[0].somModel.tcam_data[4][278][0]=80'h000000000000008f7473;
sos_loop[0].somModel.tcam_mask[4][278][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][279][0]=80'h00000000000000ff2471;
sos_loop[0].somModel.tcam_mask[4][279][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][280][0]=80'h0000000000000014b05f;
sos_loop[0].somModel.tcam_mask[4][280][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][281][0]=80'h00000000000000df9570;
sos_loop[0].somModel.tcam_mask[4][281][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][282][0]=80'h00000000000000153dbb;
sos_loop[0].somModel.tcam_mask[4][282][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][283][0]=80'h00000000000000c5d62c;
sos_loop[0].somModel.tcam_mask[4][283][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][284][0]=80'h000000000000006bf1fb;
sos_loop[0].somModel.tcam_mask[4][284][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][285][0]=80'h0000000000000025d7ea;
sos_loop[0].somModel.tcam_mask[4][285][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][286][0]=80'h000000000000007d1082;
sos_loop[0].somModel.tcam_mask[4][286][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][287][0]=80'h000000000000005f39c9;
sos_loop[0].somModel.tcam_mask[4][287][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][288][0]=80'h0000000000000009fe99;
sos_loop[0].somModel.tcam_mask[4][288][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][289][0]=80'h000000000000007b04db;
sos_loop[0].somModel.tcam_mask[4][289][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][290][0]=80'h0000000000000029dd6a;
sos_loop[0].somModel.tcam_mask[4][290][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][291][0]=80'h000000000000001fcd7e;
sos_loop[0].somModel.tcam_mask[4][291][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][292][0]=80'h000000000000005b635c;
sos_loop[0].somModel.tcam_mask[4][292][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][293][0]=80'h000000000000006eda0f;
sos_loop[0].somModel.tcam_mask[4][293][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][294][0]=80'h00000000000000cef008;
sos_loop[0].somModel.tcam_mask[4][294][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][295][0]=80'h0000000000000032dc5e;
sos_loop[0].somModel.tcam_mask[4][295][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][296][0]=80'h0000000000000050586f;
sos_loop[0].somModel.tcam_mask[4][296][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][297][0]=80'h000000000000006dc367;
sos_loop[0].somModel.tcam_mask[4][297][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][298][0]=80'h000000000000009c1de1;
sos_loop[0].somModel.tcam_mask[4][298][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][299][0]=80'h00000000000000fd77d3;
sos_loop[0].somModel.tcam_mask[4][299][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][300][0]=80'h00000000000000d3c5d4;
sos_loop[0].somModel.tcam_mask[4][300][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][301][0]=80'h000000000000000fdb0d;
sos_loop[0].somModel.tcam_mask[4][301][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][302][0]=80'h00000000000000025d51;
sos_loop[0].somModel.tcam_mask[4][302][0]=80'hfffffffffffffffc0000;
sos_loop[0].somModel.tcam_data[4][303][0]=80'h00000000000000e88800;
sos_loop[0].somModel.tcam_mask[4][303][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][304][0]=80'h00000000000000c08b8e;
sos_loop[0].somModel.tcam_mask[4][304][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][305][0]=80'h000000000000003f0392;
sos_loop[0].somModel.tcam_mask[4][305][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][306][0]=80'h00000000000000a02fb5;
sos_loop[0].somModel.tcam_mask[4][306][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][307][0]=80'h0000000000000021607f;
sos_loop[0].somModel.tcam_mask[4][307][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][308][0]=80'h000000000000008f612f;
sos_loop[0].somModel.tcam_mask[4][308][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][309][0]=80'h0000000000000034a36e;
sos_loop[0].somModel.tcam_mask[4][309][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][310][0]=80'h00000000000000899446;
sos_loop[0].somModel.tcam_mask[4][310][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][311][0]=80'h00000000000000aeaee1;
sos_loop[0].somModel.tcam_mask[4][311][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][312][0]=80'h000000000000000efa58;
sos_loop[0].somModel.tcam_mask[4][312][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][313][0]=80'h000000000000007c121d;
sos_loop[0].somModel.tcam_mask[4][313][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][314][0]=80'h0000000000000084c243;
sos_loop[0].somModel.tcam_mask[4][314][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][315][0]=80'h000000000000006fa6f1;
sos_loop[0].somModel.tcam_mask[4][315][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][316][0]=80'h00000000000000e50d93;
sos_loop[0].somModel.tcam_mask[4][316][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][317][0]=80'h0000000000000030a2f4;
sos_loop[0].somModel.tcam_mask[4][317][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][318][0]=80'h0000000000000028773f;
sos_loop[0].somModel.tcam_mask[4][318][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][319][0]=80'h000000000000000266b7;
sos_loop[0].somModel.tcam_mask[4][319][0]=80'hfffffffffffffffc0000;
sos_loop[0].somModel.tcam_data[4][320][0]=80'h00000000000000a9817d;
sos_loop[0].somModel.tcam_mask[4][320][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][321][0]=80'h000000000000003920db;
sos_loop[0].somModel.tcam_mask[4][321][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][322][0]=80'h000000000000003bfaad;
sos_loop[0].somModel.tcam_mask[4][322][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][323][0]=80'h00000000000000d9c7f1;
sos_loop[0].somModel.tcam_mask[4][323][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][324][0]=80'h000000000000005c0486;
sos_loop[0].somModel.tcam_mask[4][324][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][325][0]=80'h00000000000000d00200;
sos_loop[0].somModel.tcam_mask[4][325][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][326][0]=80'h00000000000000d49869;
sos_loop[0].somModel.tcam_mask[4][326][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][327][0]=80'h0000000000000089ee4e;
sos_loop[0].somModel.tcam_mask[4][327][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][328][0]=80'h00000000000000df942f;
sos_loop[0].somModel.tcam_mask[4][328][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][329][0]=80'h0000000000000084601d;
sos_loop[0].somModel.tcam_mask[4][329][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][330][0]=80'h000000000000001808be;
sos_loop[0].somModel.tcam_mask[4][330][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][331][0]=80'h00000000000000b502fb;
sos_loop[0].somModel.tcam_mask[4][331][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][332][0]=80'h000000000000009f2b20;
sos_loop[0].somModel.tcam_mask[4][332][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][333][0]=80'h00000000000000b2fa64;
sos_loop[0].somModel.tcam_mask[4][333][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][334][0]=80'h0000000000000080dd3b;
sos_loop[0].somModel.tcam_mask[4][334][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][335][0]=80'h0000000000000038568a;
sos_loop[0].somModel.tcam_mask[4][335][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][336][0]=80'h00000000000000ea6666;
sos_loop[0].somModel.tcam_mask[4][336][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][337][0]=80'h00000000000000dfa001;
sos_loop[0].somModel.tcam_mask[4][337][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][338][0]=80'h000000000000000396ef;
sos_loop[0].somModel.tcam_mask[4][338][0]=80'hfffffffffffffffc0000;
sos_loop[0].somModel.tcam_data[4][339][0]=80'h0000000000000061ba43;
sos_loop[0].somModel.tcam_mask[4][339][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][340][0]=80'h00000000000000080209;
sos_loop[0].somModel.tcam_mask[4][340][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][341][0]=80'h000000000000005b8fa1;
sos_loop[0].somModel.tcam_mask[4][341][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][342][0]=80'h0000000000000061c5cc;
sos_loop[0].somModel.tcam_mask[4][342][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][343][0]=80'h00000000000000b26ef1;
sos_loop[0].somModel.tcam_mask[4][343][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][344][0]=80'h00000000000000407501;
sos_loop[0].somModel.tcam_mask[4][344][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][345][0]=80'h0000000000000028ace5;
sos_loop[0].somModel.tcam_mask[4][345][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][346][0]=80'h00000000000000c579b9;
sos_loop[0].somModel.tcam_mask[4][346][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][347][0]=80'h000000000000009bfb01;
sos_loop[0].somModel.tcam_mask[4][347][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][348][0]=80'h000000000000000f34eb;
sos_loop[0].somModel.tcam_mask[4][348][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][349][0]=80'h00000000000000ab2f3d;
sos_loop[0].somModel.tcam_mask[4][349][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][350][0]=80'h00000000000000186408;
sos_loop[0].somModel.tcam_mask[4][350][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][351][0]=80'h0000000000000022a3c9;
sos_loop[0].somModel.tcam_mask[4][351][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][352][0]=80'h000000000000009aa041;
sos_loop[0].somModel.tcam_mask[4][352][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][353][0]=80'h00000000000000b46f64;
sos_loop[0].somModel.tcam_mask[4][353][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][354][0]=80'h0000000000000048548b;
sos_loop[0].somModel.tcam_mask[4][354][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][355][0]=80'h00000000000000e7ee30;
sos_loop[0].somModel.tcam_mask[4][355][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][356][0]=80'h000000000000000c7e65;
sos_loop[0].somModel.tcam_mask[4][356][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][357][0]=80'h00000000000000c4e05f;
sos_loop[0].somModel.tcam_mask[4][357][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][358][0]=80'h00000000000000cdeb94;
sos_loop[0].somModel.tcam_mask[4][358][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][359][0]=80'h00000000000000c6fbde;
sos_loop[0].somModel.tcam_mask[4][359][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][360][0]=80'h000000000000004364d2;
sos_loop[0].somModel.tcam_mask[4][360][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][361][0]=80'h0000000000000054c878;
sos_loop[0].somModel.tcam_mask[4][361][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][362][0]=80'h00000000000000244700;
sos_loop[0].somModel.tcam_mask[4][362][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][363][0]=80'h000000000000003a7f6d;
sos_loop[0].somModel.tcam_mask[4][363][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][364][0]=80'h00000000000000e03a58;
sos_loop[0].somModel.tcam_mask[4][364][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][365][0]=80'h00000000000000b0efa4;
sos_loop[0].somModel.tcam_mask[4][365][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][366][0]=80'h000000000000001e6831;
sos_loop[0].somModel.tcam_mask[4][366][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][367][0]=80'h00000000000000323acf;
sos_loop[0].somModel.tcam_mask[4][367][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][368][0]=80'h000000000000001ab23b;
sos_loop[0].somModel.tcam_mask[4][368][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][369][0]=80'h00000000000000153918;
sos_loop[0].somModel.tcam_mask[4][369][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][370][0]=80'h00000000000000a376d9;
sos_loop[0].somModel.tcam_mask[4][370][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][371][0]=80'h0000000000000066c250;
sos_loop[0].somModel.tcam_mask[4][371][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][372][0]=80'h00000000000000f46295;
sos_loop[0].somModel.tcam_mask[4][372][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][373][0]=80'h00000000000000909a33;
sos_loop[0].somModel.tcam_mask[4][373][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][374][0]=80'h00000000000000b903f6;
sos_loop[0].somModel.tcam_mask[4][374][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][375][0]=80'h00000000000000876713;
sos_loop[0].somModel.tcam_mask[4][375][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][376][0]=80'h00000000000000f203b1;
sos_loop[0].somModel.tcam_mask[4][376][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][377][0]=80'h000000000000007035e4;
sos_loop[0].somModel.tcam_mask[4][377][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][378][0]=80'h00000000000000e24033;
sos_loop[0].somModel.tcam_mask[4][378][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][379][0]=80'h00000000000000e8a4a2;
sos_loop[0].somModel.tcam_mask[4][379][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][380][0]=80'h00000000000000ece548;
sos_loop[0].somModel.tcam_mask[4][380][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][381][0]=80'h00000000000000586dfc;
sos_loop[0].somModel.tcam_mask[4][381][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][382][0]=80'h000000000000008c1319;
sos_loop[0].somModel.tcam_mask[4][382][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][383][0]=80'h00000000000000725176;
sos_loop[0].somModel.tcam_mask[4][383][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][384][0]=80'h0000000000000056cec2;
sos_loop[0].somModel.tcam_mask[4][384][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][385][0]=80'h00000000000000639a04;
sos_loop[0].somModel.tcam_mask[4][385][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][386][0]=80'h000000000000005327e0;
sos_loop[0].somModel.tcam_mask[4][386][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][387][0]=80'h000000000000001462c7;
sos_loop[0].somModel.tcam_mask[4][387][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][388][0]=80'h000000000000000d89f5;
sos_loop[0].somModel.tcam_mask[4][388][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][389][0]=80'h000000000000003902ae;
sos_loop[0].somModel.tcam_mask[4][389][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][390][0]=80'h00000000000000a2cbeb;
sos_loop[0].somModel.tcam_mask[4][390][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][391][0]=80'h000000000000000f6681;
sos_loop[0].somModel.tcam_mask[4][391][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][392][0]=80'h000000000000005dcafd;
sos_loop[0].somModel.tcam_mask[4][392][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][393][0]=80'h00000000000000691152;
sos_loop[0].somModel.tcam_mask[4][393][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][394][0]=80'h0000000000000076bcf7;
sos_loop[0].somModel.tcam_mask[4][394][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][395][0]=80'h00000000000000655333;
sos_loop[0].somModel.tcam_mask[4][395][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][396][0]=80'h0000000000000067c107;
sos_loop[0].somModel.tcam_mask[4][396][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][397][0]=80'h00000000000000bd651c;
sos_loop[0].somModel.tcam_mask[4][397][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][398][0]=80'h00000000000000d88fbe;
sos_loop[0].somModel.tcam_mask[4][398][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][399][0]=80'h000000000000003fa26a;
sos_loop[0].somModel.tcam_mask[4][399][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][400][0]=80'h00000000000000be3762;
sos_loop[0].somModel.tcam_mask[4][400][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][401][0]=80'h00000000000000ee1fc4;
sos_loop[0].somModel.tcam_mask[4][401][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][402][0]=80'h00000000000000b30bdf;
sos_loop[0].somModel.tcam_mask[4][402][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][403][0]=80'h00000000000000977fec;
sos_loop[0].somModel.tcam_mask[4][403][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][404][0]=80'h00000000000000f34eee;
sos_loop[0].somModel.tcam_mask[4][404][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][405][0]=80'h0000000000000088c78e;
sos_loop[0].somModel.tcam_mask[4][405][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][406][0]=80'h0000000000000050186a;
sos_loop[0].somModel.tcam_mask[4][406][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][407][0]=80'h0000000000000022c496;
sos_loop[0].somModel.tcam_mask[4][407][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][408][0]=80'h0000000000000074ba14;
sos_loop[0].somModel.tcam_mask[4][408][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][409][0]=80'h000000000000005fa922;
sos_loop[0].somModel.tcam_mask[4][409][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][410][0]=80'h0000000000000009f94e;
sos_loop[0].somModel.tcam_mask[4][410][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][411][0]=80'h0000000000000066d9fb;
sos_loop[0].somModel.tcam_mask[4][411][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][412][0]=80'h0000000000000010bb50;
sos_loop[0].somModel.tcam_mask[4][412][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][413][0]=80'h00000000000000139b8e;
sos_loop[0].somModel.tcam_mask[4][413][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][414][0]=80'h0000000000000034094f;
sos_loop[0].somModel.tcam_mask[4][414][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][415][0]=80'h00000000000000f852df;
sos_loop[0].somModel.tcam_mask[4][415][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][416][0]=80'h00000000000000b4b4a5;
sos_loop[0].somModel.tcam_mask[4][416][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][417][0]=80'h000000000000007de478;
sos_loop[0].somModel.tcam_mask[4][417][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][418][0]=80'h000000000000003db18f;
sos_loop[0].somModel.tcam_mask[4][418][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][419][0]=80'h00000000000000d272a2;
sos_loop[0].somModel.tcam_mask[4][419][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][420][0]=80'h000000000000008fb4b5;
sos_loop[0].somModel.tcam_mask[4][420][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][421][0]=80'h0000000000000039e1a2;
sos_loop[0].somModel.tcam_mask[4][421][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][422][0]=80'h00000000000000bcc07b;
sos_loop[0].somModel.tcam_mask[4][422][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][423][0]=80'h00000000000000b2ab05;
sos_loop[0].somModel.tcam_mask[4][423][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][424][0]=80'h00000000000000f3b478;
sos_loop[0].somModel.tcam_mask[4][424][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][425][0]=80'h000000000000009c9331;
sos_loop[0].somModel.tcam_mask[4][425][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][426][0]=80'h000000000000000570f8;
sos_loop[0].somModel.tcam_mask[4][426][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][427][0]=80'h0000000000000092489c;
sos_loop[0].somModel.tcam_mask[4][427][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][428][0]=80'h00000000000000d0fc4d;
sos_loop[0].somModel.tcam_mask[4][428][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][429][0]=80'h000000000000002acd7b;
sos_loop[0].somModel.tcam_mask[4][429][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][430][0]=80'h00000000000000ab42dd;
sos_loop[0].somModel.tcam_mask[4][430][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][431][0]=80'h00000000000000e77e1b;
sos_loop[0].somModel.tcam_mask[4][431][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][432][0]=80'h0000000000000081a3c5;
sos_loop[0].somModel.tcam_mask[4][432][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][433][0]=80'h000000000000006cf1fa;
sos_loop[0].somModel.tcam_mask[4][433][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][434][0]=80'h0000000000000034d05e;
sos_loop[0].somModel.tcam_mask[4][434][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][435][0]=80'h000000000000002b443d;
sos_loop[0].somModel.tcam_mask[4][435][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][436][0]=80'h0000000000000097d73f;
sos_loop[0].somModel.tcam_mask[4][436][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][437][0]=80'h00000000000000158478;
sos_loop[0].somModel.tcam_mask[4][437][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][438][0]=80'h00000000000000e145aa;
sos_loop[0].somModel.tcam_mask[4][438][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][439][0]=80'h000000000000001c385e;
sos_loop[0].somModel.tcam_mask[4][439][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][440][0]=80'h00000000000000adbce3;
sos_loop[0].somModel.tcam_mask[4][440][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][441][0]=80'h00000000000000d72c20;
sos_loop[0].somModel.tcam_mask[4][441][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][442][0]=80'h000000000000005a3b1b;
sos_loop[0].somModel.tcam_mask[4][442][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][443][0]=80'h000000000000005eaede;
sos_loop[0].somModel.tcam_mask[4][443][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][444][0]=80'h00000000000000651848;
sos_loop[0].somModel.tcam_mask[4][444][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][445][0]=80'h00000000000000977b39;
sos_loop[0].somModel.tcam_mask[4][445][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][446][0]=80'h000000000000005cea8e;
sos_loop[0].somModel.tcam_mask[4][446][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][447][0]=80'h000000000000003b6c9a;
sos_loop[0].somModel.tcam_mask[4][447][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][448][0]=80'h00000000000000492ee4;
sos_loop[0].somModel.tcam_mask[4][448][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][449][0]=80'h000000000000009a047c;
sos_loop[0].somModel.tcam_mask[4][449][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][450][0]=80'h00000000000000608036;
sos_loop[0].somModel.tcam_mask[4][450][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][451][0]=80'h00000000000000cbe70e;
sos_loop[0].somModel.tcam_mask[4][451][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][452][0]=80'h000000000000001eb27a;
sos_loop[0].somModel.tcam_mask[4][452][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][453][0]=80'h00000000000000751c3a;
sos_loop[0].somModel.tcam_mask[4][453][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][454][0]=80'h000000000000002b749f;
sos_loop[0].somModel.tcam_mask[4][454][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][455][0]=80'h000000000000007ab9cd;
sos_loop[0].somModel.tcam_mask[4][455][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][456][0]=80'h00000000000000db74b0;
sos_loop[0].somModel.tcam_mask[4][456][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][457][0]=80'h0000000000000038ccf5;
sos_loop[0].somModel.tcam_mask[4][457][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][458][0]=80'h00000000000000b81901;
sos_loop[0].somModel.tcam_mask[4][458][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][459][0]=80'h00000000000000db6f8a;
sos_loop[0].somModel.tcam_mask[4][459][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][460][0]=80'h00000000000000bdfaee;
sos_loop[0].somModel.tcam_mask[4][460][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][461][0]=80'h00000000000000ab9134;
sos_loop[0].somModel.tcam_mask[4][461][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][462][0]=80'h000000000000006d74aa;
sos_loop[0].somModel.tcam_mask[4][462][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][463][0]=80'h00000000000000f71076;
sos_loop[0].somModel.tcam_mask[4][463][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][464][0]=80'h00000000000000579bdc;
sos_loop[0].somModel.tcam_mask[4][464][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][465][0]=80'h00000000000000bbbd64;
sos_loop[0].somModel.tcam_mask[4][465][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][466][0]=80'h0000000000000083ae74;
sos_loop[0].somModel.tcam_mask[4][466][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][467][0]=80'h00000000000000f8c1d9;
sos_loop[0].somModel.tcam_mask[4][467][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][468][0]=80'h00000000000000c8ed3e;
sos_loop[0].somModel.tcam_mask[4][468][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][469][0]=80'h000000000000002bf8dc;
sos_loop[0].somModel.tcam_mask[4][469][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][470][0]=80'h0000000000000016e5de;
sos_loop[0].somModel.tcam_mask[4][470][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][471][0]=80'h00000000000000b99492;
sos_loop[0].somModel.tcam_mask[4][471][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][472][0]=80'h00000000000000820b16;
sos_loop[0].somModel.tcam_mask[4][472][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][473][0]=80'h000000000000008ae9cf;
sos_loop[0].somModel.tcam_mask[4][473][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][474][0]=80'h00000000000000f6aad1;
sos_loop[0].somModel.tcam_mask[4][474][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][475][0]=80'h00000000000000def433;
sos_loop[0].somModel.tcam_mask[4][475][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][476][0]=80'h0000000000000060e02b;
sos_loop[0].somModel.tcam_mask[4][476][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][477][0]=80'h00000000000000ba10d9;
sos_loop[0].somModel.tcam_mask[4][477][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][478][0]=80'h00000000000000125ae0;
sos_loop[0].somModel.tcam_mask[4][478][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][479][0]=80'h0000000000000075abca;
sos_loop[0].somModel.tcam_mask[4][479][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][480][0]=80'h000000000000007d0a37;
sos_loop[0].somModel.tcam_mask[4][480][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][481][0]=80'h0000000000000076c3eb;
sos_loop[0].somModel.tcam_mask[4][481][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][482][0]=80'h00000000000000ee5867;
sos_loop[0].somModel.tcam_mask[4][482][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][483][0]=80'h00000000000000a63aa9;
sos_loop[0].somModel.tcam_mask[4][483][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][484][0]=80'h000000000000003bf1a7;
sos_loop[0].somModel.tcam_mask[4][484][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][485][0]=80'h0000000000000041b00e;
sos_loop[0].somModel.tcam_mask[4][485][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][486][0]=80'h000000000000005dfcea;
sos_loop[0].somModel.tcam_mask[4][486][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][487][0]=80'h00000000000000856939;
sos_loop[0].somModel.tcam_mask[4][487][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][488][0]=80'h0000000000000007fdd0;
sos_loop[0].somModel.tcam_mask[4][488][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][489][0]=80'h00000000000000cac855;
sos_loop[0].somModel.tcam_mask[4][489][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][490][0]=80'h0000000000000082c86b;
sos_loop[0].somModel.tcam_mask[4][490][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][491][0]=80'h000000000000007d64e0;
sos_loop[0].somModel.tcam_mask[4][491][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][492][0]=80'h00000000000000c05790;
sos_loop[0].somModel.tcam_mask[4][492][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][493][0]=80'h0000000000000041b488;
sos_loop[0].somModel.tcam_mask[4][493][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][494][0]=80'h0000000000000019ef12;
sos_loop[0].somModel.tcam_mask[4][494][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][495][0]=80'h0000000000000089d14b;
sos_loop[0].somModel.tcam_mask[4][495][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][496][0]=80'h00000000000000b42732;
sos_loop[0].somModel.tcam_mask[4][496][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][497][0]=80'h00000000000000a795fa;
sos_loop[0].somModel.tcam_mask[4][497][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][498][0]=80'h00000000000000a72e70;
sos_loop[0].somModel.tcam_mask[4][498][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][499][0]=80'h00000000000000a16e73;
sos_loop[0].somModel.tcam_mask[4][499][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][500][0]=80'h0000000000000080fe5c;
sos_loop[0].somModel.tcam_mask[4][500][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][501][0]=80'h00000000000000bdf1f7;
sos_loop[0].somModel.tcam_mask[4][501][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][502][0]=80'h0000000000000024e03d;
sos_loop[0].somModel.tcam_mask[4][502][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][503][0]=80'h00000000000000cd8833;
sos_loop[0].somModel.tcam_mask[4][503][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][504][0]=80'h00000000000000d48427;
sos_loop[0].somModel.tcam_mask[4][504][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][505][0]=80'h0000000000000029413e;
sos_loop[0].somModel.tcam_mask[4][505][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][506][0]=80'h0000000000000099f215;
sos_loop[0].somModel.tcam_mask[4][506][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][507][0]=80'h0000000000000043ea2c;
sos_loop[0].somModel.tcam_mask[4][507][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][508][0]=80'h00000000000000b05ed6;
sos_loop[0].somModel.tcam_mask[4][508][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][509][0]=80'h00000000000000359c4e;
sos_loop[0].somModel.tcam_mask[4][509][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][510][0]=80'h00000000000000a53a50;
sos_loop[0].somModel.tcam_mask[4][510][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][511][0]=80'h00000000000000ba0217;
sos_loop[0].somModel.tcam_mask[4][511][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][512][0]=80'h00000000000000a7a8be;
sos_loop[0].somModel.tcam_mask[4][512][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][513][0]=80'h00000000000000117261;
sos_loop[0].somModel.tcam_mask[4][513][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][514][0]=80'h00000000000000ba40b1;
sos_loop[0].somModel.tcam_mask[4][514][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][515][0]=80'h00000000000000d3778c;
sos_loop[0].somModel.tcam_mask[4][515][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][516][0]=80'h00000000000000133300;
sos_loop[0].somModel.tcam_mask[4][516][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][517][0]=80'h000000000000008026d0;
sos_loop[0].somModel.tcam_mask[4][517][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][518][0]=80'h000000000000003c2a96;
sos_loop[0].somModel.tcam_mask[4][518][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][519][0]=80'h00000000000000af2172;
sos_loop[0].somModel.tcam_mask[4][519][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][520][0]=80'h00000000000000f83e69;
sos_loop[0].somModel.tcam_mask[4][520][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][521][0]=80'h000000000000002bae72;
sos_loop[0].somModel.tcam_mask[4][521][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][522][0]=80'h00000000000000aaffe3;
sos_loop[0].somModel.tcam_mask[4][522][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][523][0]=80'h00000000000000e47a3a;
sos_loop[0].somModel.tcam_mask[4][523][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][524][0]=80'h00000000000000ecf185;
sos_loop[0].somModel.tcam_mask[4][524][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][525][0]=80'h000000000000002ed0f5;
sos_loop[0].somModel.tcam_mask[4][525][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][526][0]=80'h00000000000000d53425;
sos_loop[0].somModel.tcam_mask[4][526][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][527][0]=80'h00000000000000ecfd2a;
sos_loop[0].somModel.tcam_mask[4][527][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][528][0]=80'h00000000000000c133a2;
sos_loop[0].somModel.tcam_mask[4][528][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][529][0]=80'h00000000000000b51947;
sos_loop[0].somModel.tcam_mask[4][529][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][530][0]=80'h000000000000001f5b10;
sos_loop[0].somModel.tcam_mask[4][530][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][531][0]=80'h00000000000000724175;
sos_loop[0].somModel.tcam_mask[4][531][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][532][0]=80'h000000000000004a6946;
sos_loop[0].somModel.tcam_mask[4][532][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][533][0]=80'h00000000000000f4634a;
sos_loop[0].somModel.tcam_mask[4][533][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][534][0]=80'h0000000000000074e5f6;
sos_loop[0].somModel.tcam_mask[4][534][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][535][0]=80'h00000000000000b53980;
sos_loop[0].somModel.tcam_mask[4][535][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][536][0]=80'h00000000000000bbd32a;
sos_loop[0].somModel.tcam_mask[4][536][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][537][0]=80'h000000000000004beff2;
sos_loop[0].somModel.tcam_mask[4][537][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][538][0]=80'h00000000000000c8358f;
sos_loop[0].somModel.tcam_mask[4][538][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][539][0]=80'h00000000000000cb9cd4;
sos_loop[0].somModel.tcam_mask[4][539][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][540][0]=80'h000000000000005a3371;
sos_loop[0].somModel.tcam_mask[4][540][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][541][0]=80'h00000000000000b24300;
sos_loop[0].somModel.tcam_mask[4][541][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][542][0]=80'h000000000000001fb996;
sos_loop[0].somModel.tcam_mask[4][542][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][543][0]=80'h00000000000000bd4f61;
sos_loop[0].somModel.tcam_mask[4][543][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][544][0]=80'h000000000000008abbcd;
sos_loop[0].somModel.tcam_mask[4][544][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][545][0]=80'h00000000000000b9b2c6;
sos_loop[0].somModel.tcam_mask[4][545][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][546][0]=80'h00000000000000638408;
sos_loop[0].somModel.tcam_mask[4][546][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][547][0]=80'h00000000000000d821e0;
sos_loop[0].somModel.tcam_mask[4][547][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][548][0]=80'h00000000000000694d89;
sos_loop[0].somModel.tcam_mask[4][548][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][549][0]=80'h00000000000000cc2430;
sos_loop[0].somModel.tcam_mask[4][549][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][550][0]=80'h000000000000000b3c95;
sos_loop[0].somModel.tcam_mask[4][550][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][551][0]=80'h000000000000002c40c9;
sos_loop[0].somModel.tcam_mask[4][551][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][552][0]=80'h00000000000000ec7053;
sos_loop[0].somModel.tcam_mask[4][552][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][553][0]=80'h000000000000008adfbd;
sos_loop[0].somModel.tcam_mask[4][553][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][554][0]=80'h0000000000000015e421;
sos_loop[0].somModel.tcam_mask[4][554][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][555][0]=80'h00000000000000cd639d;
sos_loop[0].somModel.tcam_mask[4][555][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][556][0]=80'h0000000000000006a5ec;
sos_loop[0].somModel.tcam_mask[4][556][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][557][0]=80'h000000000000004837b3;
sos_loop[0].somModel.tcam_mask[4][557][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][558][0]=80'h000000000000003c1296;
sos_loop[0].somModel.tcam_mask[4][558][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][559][0]=80'h000000000000009854db;
sos_loop[0].somModel.tcam_mask[4][559][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][560][0]=80'h00000000000000e23953;
sos_loop[0].somModel.tcam_mask[4][560][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][561][0]=80'h000000000000006e5f61;
sos_loop[0].somModel.tcam_mask[4][561][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][562][0]=80'h00000000000000b67704;
sos_loop[0].somModel.tcam_mask[4][562][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][563][0]=80'h00000000000000c188f5;
sos_loop[0].somModel.tcam_mask[4][563][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][564][0]=80'h000000000000009f0af0;
sos_loop[0].somModel.tcam_mask[4][564][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][565][0]=80'h0000000000000013deba;
sos_loop[0].somModel.tcam_mask[4][565][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][566][0]=80'h00000000000000d836a2;
sos_loop[0].somModel.tcam_mask[4][566][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][567][0]=80'h00000000000000378015;
sos_loop[0].somModel.tcam_mask[4][567][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][568][0]=80'h0000000000000006857c;
sos_loop[0].somModel.tcam_mask[4][568][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][569][0]=80'h00000000000000920848;
sos_loop[0].somModel.tcam_mask[4][569][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][570][0]=80'h00000000000000df91e5;
sos_loop[0].somModel.tcam_mask[4][570][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][571][0]=80'h00000000000000203539;
sos_loop[0].somModel.tcam_mask[4][571][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][572][0]=80'h00000000000000e0e16e;
sos_loop[0].somModel.tcam_mask[4][572][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][573][0]=80'h00000000000000518348;
sos_loop[0].somModel.tcam_mask[4][573][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][574][0]=80'h0000000000000029589f;
sos_loop[0].somModel.tcam_mask[4][574][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][575][0]=80'h00000000000000d5eff5;
sos_loop[0].somModel.tcam_mask[4][575][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][576][0]=80'h00000000000000a8909a;
sos_loop[0].somModel.tcam_mask[4][576][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][577][0]=80'h00000000000000c6ccb7;
sos_loop[0].somModel.tcam_mask[4][577][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][578][0]=80'h000000000000008fd56d;
sos_loop[0].somModel.tcam_mask[4][578][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][579][0]=80'h00000000000000bf7f6d;
sos_loop[0].somModel.tcam_mask[4][579][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][580][0]=80'h000000000000006a229b;
sos_loop[0].somModel.tcam_mask[4][580][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][581][0]=80'h00000000000000a7dd84;
sos_loop[0].somModel.tcam_mask[4][581][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][582][0]=80'h000000000000003d9854;
sos_loop[0].somModel.tcam_mask[4][582][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][583][0]=80'h000000000000003c87c6;
sos_loop[0].somModel.tcam_mask[4][583][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][584][0]=80'h00000000000000588ad5;
sos_loop[0].somModel.tcam_mask[4][584][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][585][0]=80'h00000000000000eaaf14;
sos_loop[0].somModel.tcam_mask[4][585][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][586][0]=80'h00000000000000344bf2;
sos_loop[0].somModel.tcam_mask[4][586][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][587][0]=80'h000000000000003d9161;
sos_loop[0].somModel.tcam_mask[4][587][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][588][0]=80'h000000000000000415ce;
sos_loop[0].somModel.tcam_mask[4][588][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][589][0]=80'h000000000000000b69cc;
sos_loop[0].somModel.tcam_mask[4][589][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][590][0]=80'h00000000000000fe9312;
sos_loop[0].somModel.tcam_mask[4][590][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][591][0]=80'h00000000000000878cb6;
sos_loop[0].somModel.tcam_mask[4][591][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][592][0]=80'h0000000000000038cf4e;
sos_loop[0].somModel.tcam_mask[4][592][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][593][0]=80'h0000000000000076dcb4;
sos_loop[0].somModel.tcam_mask[4][593][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][594][0]=80'h00000000000000702f85;
sos_loop[0].somModel.tcam_mask[4][594][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][595][0]=80'h00000000000000ecdc20;
sos_loop[0].somModel.tcam_mask[4][595][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][596][0]=80'h00000000000000064eed;
sos_loop[0].somModel.tcam_mask[4][596][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][597][0]=80'h00000000000000197ad7;
sos_loop[0].somModel.tcam_mask[4][597][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][598][0]=80'h00000000000000860fe2;
sos_loop[0].somModel.tcam_mask[4][598][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][599][0]=80'h00000000000000aafcfa;
sos_loop[0].somModel.tcam_mask[4][599][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][600][0]=80'h00000000000000b3fdf0;
sos_loop[0].somModel.tcam_mask[4][600][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][601][0]=80'h00000000000000075513;
sos_loop[0].somModel.tcam_mask[4][601][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][602][0]=80'h0000000000000013141b;
sos_loop[0].somModel.tcam_mask[4][602][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][603][0]=80'h00000000000000d07c80;
sos_loop[0].somModel.tcam_mask[4][603][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][604][0]=80'h000000000000007023d5;
sos_loop[0].somModel.tcam_mask[4][604][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][605][0]=80'h0000000000000088bbc7;
sos_loop[0].somModel.tcam_mask[4][605][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][606][0]=80'h000000000000008bd1c2;
sos_loop[0].somModel.tcam_mask[4][606][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][607][0]=80'h00000000000000ede0cc;
sos_loop[0].somModel.tcam_mask[4][607][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][608][0]=80'h0000000000000011d1b8;
sos_loop[0].somModel.tcam_mask[4][608][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][609][0]=80'h00000000000000d0feb3;
sos_loop[0].somModel.tcam_mask[4][609][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][610][0]=80'h00000000000000ef7aab;
sos_loop[0].somModel.tcam_mask[4][610][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][611][0]=80'h00000000000000929846;
sos_loop[0].somModel.tcam_mask[4][611][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][612][0]=80'h0000000000000087f8f5;
sos_loop[0].somModel.tcam_mask[4][612][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][613][0]=80'h00000000000000f6d906;
sos_loop[0].somModel.tcam_mask[4][613][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][614][0]=80'h00000000000000301023;
sos_loop[0].somModel.tcam_mask[4][614][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][615][0]=80'h00000000000000c0367e;
sos_loop[0].somModel.tcam_mask[4][615][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][616][0]=80'h000000000000000b5225;
sos_loop[0].somModel.tcam_mask[4][616][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][617][0]=80'h000000000000001abda8;
sos_loop[0].somModel.tcam_mask[4][617][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][618][0]=80'h00000000000000f76cf7;
sos_loop[0].somModel.tcam_mask[4][618][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][619][0]=80'h00000000000000715672;
sos_loop[0].somModel.tcam_mask[4][619][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][620][0]=80'h000000000000007a6132;
sos_loop[0].somModel.tcam_mask[4][620][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][621][0]=80'h00000000000000443d93;
sos_loop[0].somModel.tcam_mask[4][621][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][622][0]=80'h00000000000000eb213b;
sos_loop[0].somModel.tcam_mask[4][622][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][623][0]=80'h000000000000004d47a0;
sos_loop[0].somModel.tcam_mask[4][623][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][624][0]=80'h00000000000000a05377;
sos_loop[0].somModel.tcam_mask[4][624][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][625][0]=80'h000000000000006ac1b8;
sos_loop[0].somModel.tcam_mask[4][625][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][626][0]=80'h000000000000007a773d;
sos_loop[0].somModel.tcam_mask[4][626][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][627][0]=80'h00000000000000e5e3a5;
sos_loop[0].somModel.tcam_mask[4][627][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][628][0]=80'h00000000000000c9746b;
sos_loop[0].somModel.tcam_mask[4][628][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][629][0]=80'h0000000000000023a9d3;
sos_loop[0].somModel.tcam_mask[4][629][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][630][0]=80'h000000000000004ec356;
sos_loop[0].somModel.tcam_mask[4][630][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][631][0]=80'h00000000000000075d68;
sos_loop[0].somModel.tcam_mask[4][631][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][632][0]=80'h000000000000003f8eba;
sos_loop[0].somModel.tcam_mask[4][632][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][633][0]=80'h000000000000004d98e8;
sos_loop[0].somModel.tcam_mask[4][633][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][634][0]=80'h0000000000000098da92;
sos_loop[0].somModel.tcam_mask[4][634][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][635][0]=80'h00000000000000ca02ef;
sos_loop[0].somModel.tcam_mask[4][635][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][636][0]=80'h00000000000000924656;
sos_loop[0].somModel.tcam_mask[4][636][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][637][0]=80'h000000000000004eb306;
sos_loop[0].somModel.tcam_mask[4][637][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][638][0]=80'h0000000000000033a608;
sos_loop[0].somModel.tcam_mask[4][638][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][639][0]=80'h00000000000000291e21;
sos_loop[0].somModel.tcam_mask[4][639][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][640][0]=80'h00000000000000c4dc56;
sos_loop[0].somModel.tcam_mask[4][640][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][641][0]=80'h000000000000001b53a4;
sos_loop[0].somModel.tcam_mask[4][641][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][642][0]=80'h0000000000000009d22f;
sos_loop[0].somModel.tcam_mask[4][642][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][643][0]=80'h000000000000005a1b8f;
sos_loop[0].somModel.tcam_mask[4][643][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][644][0]=80'h00000000000000e01679;
sos_loop[0].somModel.tcam_mask[4][644][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][645][0]=80'h0000000000000044e0ed;
sos_loop[0].somModel.tcam_mask[4][645][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][646][0]=80'h00000000000000c9bb74;
sos_loop[0].somModel.tcam_mask[4][646][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][647][0]=80'h000000000000005c1683;
sos_loop[0].somModel.tcam_mask[4][647][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][648][0]=80'h000000000000005fbc9d;
sos_loop[0].somModel.tcam_mask[4][648][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][649][0]=80'h00000000000000bc2b03;
sos_loop[0].somModel.tcam_mask[4][649][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][650][0]=80'h0000000000000044df86;
sos_loop[0].somModel.tcam_mask[4][650][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][651][0]=80'h00000000000000dadec5;
sos_loop[0].somModel.tcam_mask[4][651][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][652][0]=80'h000000000000002fa3c2;
sos_loop[0].somModel.tcam_mask[4][652][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][653][0]=80'h00000000000000795c0b;
sos_loop[0].somModel.tcam_mask[4][653][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][654][0]=80'h00000000000000c6f84e;
sos_loop[0].somModel.tcam_mask[4][654][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][655][0]=80'h00000000000000b16934;
sos_loop[0].somModel.tcam_mask[4][655][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][656][0]=80'h000000000000009460ec;
sos_loop[0].somModel.tcam_mask[4][656][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][657][0]=80'h00000000000000961e88;
sos_loop[0].somModel.tcam_mask[4][657][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][658][0]=80'h00000000000000c93603;
sos_loop[0].somModel.tcam_mask[4][658][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][659][0]=80'h00000000000000f71bb0;
sos_loop[0].somModel.tcam_mask[4][659][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][660][0]=80'h00000000000000b1611c;
sos_loop[0].somModel.tcam_mask[4][660][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][661][0]=80'h00000000000000ec7932;
sos_loop[0].somModel.tcam_mask[4][661][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][662][0]=80'h0000000000000043bb09;
sos_loop[0].somModel.tcam_mask[4][662][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][663][0]=80'h00000000000000040cb8;
sos_loop[0].somModel.tcam_mask[4][663][0]=80'hfffffffffffffff80000;
sos_loop[0].somModel.tcam_data[4][664][0]=80'h0000000000000085d475;
sos_loop[0].somModel.tcam_mask[4][664][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][665][0]=80'h00000000000000a661a8;
sos_loop[0].somModel.tcam_mask[4][665][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][666][0]=80'h000000000000000f38b5;
sos_loop[0].somModel.tcam_mask[4][666][0]=80'hfffffffffffffff00000;
sos_loop[0].somModel.tcam_data[4][667][0]=80'h00000000000000986622;
sos_loop[0].somModel.tcam_mask[4][667][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][668][0]=80'h0000000000000072876e;
sos_loop[0].somModel.tcam_mask[4][668][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][669][0]=80'h0000000000000026c981;
sos_loop[0].somModel.tcam_mask[4][669][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][670][0]=80'h00000000000000c3c23a;
sos_loop[0].somModel.tcam_mask[4][670][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][671][0]=80'h00000000000000907259;
sos_loop[0].somModel.tcam_mask[4][671][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][672][0]=80'h0000000000000052165d;
sos_loop[0].somModel.tcam_mask[4][672][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][673][0]=80'h0000000000000095fcd7;
sos_loop[0].somModel.tcam_mask[4][673][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][674][0]=80'h000000000000002dc5de;
sos_loop[0].somModel.tcam_mask[4][674][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][675][0]=80'h000000000000003bd5a3;
sos_loop[0].somModel.tcam_mask[4][675][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][676][0]=80'h00000000000000a551ba;
sos_loop[0].somModel.tcam_mask[4][676][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][677][0]=80'h0000000000000035e5cb;
sos_loop[0].somModel.tcam_mask[4][677][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][678][0]=80'h00000000000000c960bd;
sos_loop[0].somModel.tcam_mask[4][678][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][679][0]=80'h0000000000000023b8b6;
sos_loop[0].somModel.tcam_mask[4][679][0]=80'hffffffffffffffc00000;
sos_loop[0].somModel.tcam_data[4][680][0]=80'h00000000000000d4d778;
sos_loop[0].somModel.tcam_mask[4][680][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][681][0]=80'h00000000000000ea3ee3;
sos_loop[0].somModel.tcam_mask[4][681][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][682][0]=80'h000000000000001d84d3;
sos_loop[0].somModel.tcam_mask[4][682][0]=80'hffffffffffffffe00000;
sos_loop[0].somModel.tcam_data[4][683][0]=80'h0000000000000077135c;
sos_loop[0].somModel.tcam_mask[4][683][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][684][0]=80'h0000000000000061df00;
sos_loop[0].somModel.tcam_mask[4][684][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][685][0]=80'h00000000000000a9a5bc;
sos_loop[0].somModel.tcam_mask[4][685][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][686][0]=80'h00000000000000ba4d19;
sos_loop[0].somModel.tcam_mask[4][686][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][687][0]=80'h00000000000000ccf409;
sos_loop[0].somModel.tcam_mask[4][687][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][688][0]=80'h0000000000000085da8d;
sos_loop[0].somModel.tcam_mask[4][688][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][689][0]=80'h00000000000000615d80;
sos_loop[0].somModel.tcam_mask[4][689][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][690][0]=80'h00000000000000726469;
sos_loop[0].somModel.tcam_mask[4][690][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][691][0]=80'h0000000000000069cc0a;
sos_loop[0].somModel.tcam_mask[4][691][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][692][0]=80'h00000000000000b23db7;
sos_loop[0].somModel.tcam_mask[4][692][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][693][0]=80'h00000000000000512c45;
sos_loop[0].somModel.tcam_mask[4][693][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][694][0]=80'h00000000000000dcffc3;
sos_loop[0].somModel.tcam_mask[4][694][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][695][0]=80'h00000000000000cc8fd4;
sos_loop[0].somModel.tcam_mask[4][695][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][696][0]=80'h00000000000000ac910e;
sos_loop[0].somModel.tcam_mask[4][696][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][697][0]=80'h0000000000000066efed;
sos_loop[0].somModel.tcam_mask[4][697][0]=80'hffffffffffffff800000;
sos_loop[0].somModel.tcam_data[4][698][0]=80'h00000000000000d0094e;
sos_loop[0].somModel.tcam_mask[4][698][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][699][0]=80'h00000000000000c23370;
sos_loop[0].somModel.tcam_mask[4][699][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.tcam_data[4][700][0]=80'h00000000000000ace597;
sos_loop[0].somModel.tcam_mask[4][700][0]=80'hffffffffffffff000000;
sos_loop[0].somModel.sram_dat[4][0][0]=96'hdeadbf;
sos_loop[0].somModel.sram_ptr[4][0]=939;
sos_loop[0].somModel.sram_dat[4][1][0]=96'h5b391854;
sos_loop[0].somModel.sram_ptr[4][1]=3;
sos_loop[0].somModel.sram_dat[4][2][0]=96'h3e47f882;
sos_loop[0].somModel.sram_ptr[4][2]=3;
sos_loop[0].somModel.sram_dat[4][3][0]=96'h5914e02b;
sos_loop[0].somModel.sram_ptr[4][3]=3;
sos_loop[0].somModel.sram_dat[4][4][0]=96'h4195b117;
sos_loop[0].somModel.sram_ptr[4][4]=3;
sos_loop[0].somModel.sram_dat[4][5][0]=96'h66a71524;
sos_loop[0].somModel.sram_ptr[4][5]=3;
sos_loop[0].somModel.sram_dat[4][6][0]=96'h51451b67;
sos_loop[0].somModel.sram_ptr[4][6]=3;
sos_loop[0].somModel.sram_dat[4][7][0]=96'h21189ffb;
sos_loop[0].somModel.sram_ptr[4][7]=3;
sos_loop[0].somModel.sram_dat[4][8][0]=96'hcbc0b312;
sos_loop[0].somModel.sram_ptr[4][8]=3;
sos_loop[0].somModel.sram_dat[4][9][0]=96'h2d22c053;
sos_loop[0].somModel.sram_ptr[4][9]=3;
sos_loop[0].somModel.sram_dat[4][10][0]=96'hb3cdad1c;
sos_loop[0].somModel.sram_ptr[4][10]=3;
sos_loop[0].somModel.sram_dat[4][11][0]=96'hf1426fee;
sos_loop[0].somModel.sram_ptr[4][11]=3;
sos_loop[0].somModel.sram_dat[4][12][0]=96'h58f695e9;
sos_loop[0].somModel.sram_ptr[4][12]=3;
sos_loop[0].somModel.sram_dat[4][13][0]=96'h8c8a5f2f;
sos_loop[0].somModel.sram_ptr[4][13]=3;
sos_loop[0].somModel.sram_dat[4][14][0]=96'ha4687d04;
sos_loop[0].somModel.sram_ptr[4][14]=3;
sos_loop[0].somModel.sram_dat[4][15][0]=96'hcda417ee;
sos_loop[0].somModel.sram_ptr[4][15]=3;
sos_loop[0].somModel.sram_dat[4][16][0]=96'hcc1a14c9;
sos_loop[0].somModel.sram_ptr[4][16]=3;
sos_loop[0].somModel.sram_dat[4][17][0]=96'hda52651a;
sos_loop[0].somModel.sram_ptr[4][17]=3;
sos_loop[0].somModel.sram_dat[4][18][0]=96'h86df7509;
sos_loop[0].somModel.sram_ptr[4][18]=3;
sos_loop[0].somModel.sram_dat[4][19][0]=96'h4d81cf6e;
sos_loop[0].somModel.sram_ptr[4][19]=3;
sos_loop[0].somModel.sram_dat[4][20][0]=96'hbbe63f40;
sos_loop[0].somModel.sram_ptr[4][20]=3;
sos_loop[0].somModel.sram_dat[4][21][0]=96'ha2d47841;
sos_loop[0].somModel.sram_ptr[4][21]=3;
sos_loop[0].somModel.sram_dat[4][22][0]=96'h24aa1d23;
sos_loop[0].somModel.sram_ptr[4][22]=3;
sos_loop[0].somModel.sram_dat[4][23][0]=96'h83a28630;
sos_loop[0].somModel.sram_ptr[4][23]=3;
sos_loop[0].somModel.sram_dat[4][24][0]=96'hf752362;
sos_loop[0].somModel.sram_ptr[4][24]=3;
sos_loop[0].somModel.sram_dat[4][25][0]=96'hcf1da1db;
sos_loop[0].somModel.sram_ptr[4][25]=3;
sos_loop[0].somModel.sram_dat[4][26][0]=96'h5355e83;
sos_loop[0].somModel.sram_ptr[4][26]=3;
sos_loop[0].somModel.sram_dat[4][27][0]=96'hb96a09bb;
sos_loop[0].somModel.sram_ptr[4][27]=3;
sos_loop[0].somModel.sram_dat[4][28][0]=96'hc02936d5;
sos_loop[0].somModel.sram_ptr[4][28]=3;
sos_loop[0].somModel.sram_dat[4][29][0]=96'h5d6d63e1;
sos_loop[0].somModel.sram_ptr[4][29]=3;
sos_loop[0].somModel.sram_dat[4][30][0]=96'hfbf7c266;
sos_loop[0].somModel.sram_ptr[4][30]=3;
sos_loop[0].somModel.sram_dat[4][31][0]=96'hb357e4e5;
sos_loop[0].somModel.sram_ptr[4][31]=3;
sos_loop[0].somModel.sram_dat[4][32][0]=96'h9b1fb39b;
sos_loop[0].somModel.sram_ptr[4][32]=3;
sos_loop[0].somModel.sram_dat[4][33][0]=96'h52fb9bde;
sos_loop[0].somModel.sram_ptr[4][33]=3;
sos_loop[0].somModel.sram_dat[4][34][0]=96'hfca1984d;
sos_loop[0].somModel.sram_ptr[4][34]=3;
sos_loop[0].somModel.sram_dat[4][35][0]=96'h740649d4;
sos_loop[0].somModel.sram_ptr[4][35]=3;
sos_loop[0].somModel.sram_dat[4][36][0]=96'h9fe5838f;
sos_loop[0].somModel.sram_ptr[4][36]=3;
sos_loop[0].somModel.sram_dat[4][37][0]=96'hd0e352d5;
sos_loop[0].somModel.sram_ptr[4][37]=3;
sos_loop[0].somModel.sram_dat[4][38][0]=96'hec62b4dc;
sos_loop[0].somModel.sram_ptr[4][38]=3;
sos_loop[0].somModel.sram_dat[4][39][0]=96'hc36e613b;
sos_loop[0].somModel.sram_ptr[4][39]=3;
sos_loop[0].somModel.sram_dat[4][40][0]=96'h5479fe;
sos_loop[0].somModel.sram_ptr[4][40]=3;
sos_loop[0].somModel.sram_dat[4][41][0]=96'hdbd26ba9;
sos_loop[0].somModel.sram_ptr[4][41]=3;
sos_loop[0].somModel.sram_dat[4][42][0]=96'hd6df9413;
sos_loop[0].somModel.sram_ptr[4][42]=3;
sos_loop[0].somModel.sram_dat[4][43][0]=96'hc385e52b;
sos_loop[0].somModel.sram_ptr[4][43]=3;
sos_loop[0].somModel.sram_dat[4][44][0]=96'hc476407e;
sos_loop[0].somModel.sram_ptr[4][44]=3;
sos_loop[0].somModel.sram_dat[4][45][0]=96'h25bb9adf;
sos_loop[0].somModel.sram_ptr[4][45]=3;
sos_loop[0].somModel.sram_dat[4][46][0]=96'hafef0d47;
sos_loop[0].somModel.sram_ptr[4][46]=3;
sos_loop[0].somModel.sram_dat[4][47][0]=96'h1b798fdf;
sos_loop[0].somModel.sram_ptr[4][47]=3;
sos_loop[0].somModel.sram_dat[4][48][0]=96'h31a3da4a;
sos_loop[0].somModel.sram_ptr[4][48]=3;
sos_loop[0].somModel.sram_dat[4][49][0]=96'hc5ed41ab;
sos_loop[0].somModel.sram_ptr[4][49]=3;
sos_loop[0].somModel.sram_dat[4][50][0]=96'hba3cc864;
sos_loop[0].somModel.sram_ptr[4][50]=3;
sos_loop[0].somModel.sram_dat[4][51][0]=96'h32ef62f2;
sos_loop[0].somModel.sram_ptr[4][51]=3;
sos_loop[0].somModel.sram_dat[4][52][0]=96'h6c4301a5;
sos_loop[0].somModel.sram_ptr[4][52]=3;
sos_loop[0].somModel.sram_dat[4][53][0]=96'h235a7415;
sos_loop[0].somModel.sram_ptr[4][53]=3;
sos_loop[0].somModel.sram_dat[4][54][0]=96'he83475e2;
sos_loop[0].somModel.sram_ptr[4][54]=3;
sos_loop[0].somModel.sram_dat[4][55][0]=96'h5efe85e6;
sos_loop[0].somModel.sram_ptr[4][55]=3;
sos_loop[0].somModel.sram_dat[4][56][0]=96'hbb4b49f8;
sos_loop[0].somModel.sram_ptr[4][56]=3;
sos_loop[0].somModel.sram_dat[4][57][0]=96'hdf9df74d;
sos_loop[0].somModel.sram_ptr[4][57]=3;
sos_loop[0].somModel.sram_dat[4][58][0]=96'h6633fdf5;
sos_loop[0].somModel.sram_ptr[4][58]=3;
sos_loop[0].somModel.sram_dat[4][59][0]=96'h271dda58;
sos_loop[0].somModel.sram_ptr[4][59]=3;
sos_loop[0].somModel.sram_dat[4][60][0]=96'h3b9537e2;
sos_loop[0].somModel.sram_ptr[4][60]=3;
sos_loop[0].somModel.sram_dat[4][61][0]=96'h29f59cc;
sos_loop[0].somModel.sram_ptr[4][61]=3;
sos_loop[0].somModel.sram_dat[4][62][0]=96'h214f6a30;
sos_loop[0].somModel.sram_ptr[4][62]=3;
sos_loop[0].somModel.sram_dat[4][63][0]=96'h301509db;
sos_loop[0].somModel.sram_ptr[4][63]=3;
sos_loop[0].somModel.sram_dat[4][64][0]=96'h9675af7b;
sos_loop[0].somModel.sram_ptr[4][64]=3;
sos_loop[0].somModel.sram_dat[4][65][0]=96'h623a5d56;
sos_loop[0].somModel.sram_ptr[4][65]=3;
sos_loop[0].somModel.sram_dat[4][66][0]=96'hb072e20e;
sos_loop[0].somModel.sram_ptr[4][66]=3;
sos_loop[0].somModel.sram_dat[4][67][0]=96'hff1ffbde;
sos_loop[0].somModel.sram_ptr[4][67]=3;
sos_loop[0].somModel.sram_dat[4][68][0]=96'he73e0b0f;
sos_loop[0].somModel.sram_ptr[4][68]=3;
sos_loop[0].somModel.sram_dat[4][69][0]=96'h142ef689;
sos_loop[0].somModel.sram_ptr[4][69]=3;
sos_loop[0].somModel.sram_dat[4][70][0]=96'hf1aaddea;
sos_loop[0].somModel.sram_ptr[4][70]=3;
sos_loop[0].somModel.sram_dat[4][71][0]=96'h52626454;
sos_loop[0].somModel.sram_ptr[4][71]=3;
sos_loop[0].somModel.sram_dat[4][72][0]=96'ha731740c;
sos_loop[0].somModel.sram_ptr[4][72]=3;
sos_loop[0].somModel.sram_dat[4][73][0]=96'h91de6f55;
sos_loop[0].somModel.sram_ptr[4][73]=3;
sos_loop[0].somModel.sram_dat[4][74][0]=96'h3ae6fcaa;
sos_loop[0].somModel.sram_ptr[4][74]=3;
sos_loop[0].somModel.sram_dat[4][75][0]=96'h6d454300;
sos_loop[0].somModel.sram_ptr[4][75]=3;
sos_loop[0].somModel.sram_dat[4][76][0]=96'h44403806;
sos_loop[0].somModel.sram_ptr[4][76]=3;
sos_loop[0].somModel.sram_dat[4][77][0]=96'h90a17056;
sos_loop[0].somModel.sram_ptr[4][77]=3;
sos_loop[0].somModel.sram_dat[4][78][0]=96'hd6246cf5;
sos_loop[0].somModel.sram_ptr[4][78]=3;
sos_loop[0].somModel.sram_dat[4][79][0]=96'h72c15812;
sos_loop[0].somModel.sram_ptr[4][79]=3;
sos_loop[0].somModel.sram_dat[4][80][0]=96'h9eac0e5d;
sos_loop[0].somModel.sram_ptr[4][80]=3;
sos_loop[0].somModel.sram_dat[4][81][0]=96'ha78d57a7;
sos_loop[0].somModel.sram_ptr[4][81]=3;
sos_loop[0].somModel.sram_dat[4][82][0]=96'hb5fb3b40;
sos_loop[0].somModel.sram_ptr[4][82]=3;
sos_loop[0].somModel.sram_dat[4][83][0]=96'hc6d29d2b;
sos_loop[0].somModel.sram_ptr[4][83]=3;
sos_loop[0].somModel.sram_dat[4][84][0]=96'he2e8b161;
sos_loop[0].somModel.sram_ptr[4][84]=3;
sos_loop[0].somModel.sram_dat[4][85][0]=96'hc9794b3d;
sos_loop[0].somModel.sram_ptr[4][85]=3;
sos_loop[0].somModel.sram_dat[4][86][0]=96'h662da1a8;
sos_loop[0].somModel.sram_ptr[4][86]=3;
sos_loop[0].somModel.sram_dat[4][87][0]=96'h6642c62e;
sos_loop[0].somModel.sram_ptr[4][87]=3;
sos_loop[0].somModel.sram_dat[4][88][0]=96'ha3b6c0c1;
sos_loop[0].somModel.sram_ptr[4][88]=3;
sos_loop[0].somModel.sram_dat[4][89][0]=96'hc24d613d;
sos_loop[0].somModel.sram_ptr[4][89]=3;
sos_loop[0].somModel.sram_dat[4][90][0]=96'h910917bf;
sos_loop[0].somModel.sram_ptr[4][90]=3;
sos_loop[0].somModel.sram_dat[4][91][0]=96'h3155f993;
sos_loop[0].somModel.sram_ptr[4][91]=3;
sos_loop[0].somModel.sram_dat[4][92][0]=96'h2a6f131a;
sos_loop[0].somModel.sram_ptr[4][92]=3;
sos_loop[0].somModel.sram_dat[4][93][0]=96'he3b4b767;
sos_loop[0].somModel.sram_ptr[4][93]=3;
sos_loop[0].somModel.sram_dat[4][94][0]=96'he0ae5572;
sos_loop[0].somModel.sram_ptr[4][94]=3;
sos_loop[0].somModel.sram_dat[4][95][0]=96'ha94d69c6;
sos_loop[0].somModel.sram_ptr[4][95]=3;
sos_loop[0].somModel.sram_dat[4][96][0]=96'h6195fa59;
sos_loop[0].somModel.sram_ptr[4][96]=3;
sos_loop[0].somModel.sram_dat[4][97][0]=96'h95f69846;
sos_loop[0].somModel.sram_ptr[4][97]=3;
sos_loop[0].somModel.sram_dat[4][98][0]=96'he827b8be;
sos_loop[0].somModel.sram_ptr[4][98]=3;
sos_loop[0].somModel.sram_dat[4][99][0]=96'hb8ac9596;
sos_loop[0].somModel.sram_ptr[4][99]=3;
sos_loop[0].somModel.sram_dat[4][100][0]=96'hddf142e;
sos_loop[0].somModel.sram_ptr[4][100]=3;
sos_loop[0].somModel.sram_dat[4][101][0]=96'h5314b7fd;
sos_loop[0].somModel.sram_ptr[4][101]=3;
sos_loop[0].somModel.sram_dat[4][102][0]=96'h7ea588c1;
sos_loop[0].somModel.sram_ptr[4][102]=3;
sos_loop[0].somModel.sram_dat[4][103][0]=96'haf21ab63;
sos_loop[0].somModel.sram_ptr[4][103]=3;
sos_loop[0].somModel.sram_dat[4][104][0]=96'h5eb7a1ad;
sos_loop[0].somModel.sram_ptr[4][104]=3;
sos_loop[0].somModel.sram_dat[4][105][0]=96'hdccbcdaa;
sos_loop[0].somModel.sram_ptr[4][105]=3;
sos_loop[0].somModel.sram_dat[4][106][0]=96'h626ccf1e;
sos_loop[0].somModel.sram_ptr[4][106]=3;
sos_loop[0].somModel.sram_dat[4][107][0]=96'h46c8d7ad;
sos_loop[0].somModel.sram_ptr[4][107]=3;
sos_loop[0].somModel.sram_dat[4][108][0]=96'hb278cf5a;
sos_loop[0].somModel.sram_ptr[4][108]=3;
sos_loop[0].somModel.sram_dat[4][109][0]=96'he34af42a;
sos_loop[0].somModel.sram_ptr[4][109]=3;
sos_loop[0].somModel.sram_dat[4][110][0]=96'hc927dedb;
sos_loop[0].somModel.sram_ptr[4][110]=3;
sos_loop[0].somModel.sram_dat[4][111][0]=96'hee6dd01c;
sos_loop[0].somModel.sram_ptr[4][111]=3;
sos_loop[0].somModel.sram_dat[4][112][0]=96'hdf79afea;
sos_loop[0].somModel.sram_ptr[4][112]=3;
sos_loop[0].somModel.sram_dat[4][113][0]=96'hb711e4ad;
sos_loop[0].somModel.sram_ptr[4][113]=3;
sos_loop[0].somModel.sram_dat[4][114][0]=96'h525533c2;
sos_loop[0].somModel.sram_ptr[4][114]=3;
sos_loop[0].somModel.sram_dat[4][115][0]=96'hbdc263d3;
sos_loop[0].somModel.sram_ptr[4][115]=3;
sos_loop[0].somModel.sram_dat[4][116][0]=96'h592e4945;
sos_loop[0].somModel.sram_ptr[4][116]=3;
sos_loop[0].somModel.sram_dat[4][117][0]=96'he9b90599;
sos_loop[0].somModel.sram_ptr[4][117]=3;
sos_loop[0].somModel.sram_dat[4][118][0]=96'h956729f4;
sos_loop[0].somModel.sram_ptr[4][118]=3;
sos_loop[0].somModel.sram_dat[4][119][0]=96'hf35f3a5e;
sos_loop[0].somModel.sram_ptr[4][119]=3;
sos_loop[0].somModel.sram_dat[4][120][0]=96'h7ab0f7bc;
sos_loop[0].somModel.sram_ptr[4][120]=3;
sos_loop[0].somModel.sram_dat[4][121][0]=96'h638321a1;
sos_loop[0].somModel.sram_ptr[4][121]=3;
sos_loop[0].somModel.sram_dat[4][122][0]=96'h28e8ce21;
sos_loop[0].somModel.sram_ptr[4][122]=3;
sos_loop[0].somModel.sram_dat[4][123][0]=96'h58309313;
sos_loop[0].somModel.sram_ptr[4][123]=3;
sos_loop[0].somModel.sram_dat[4][124][0]=96'h14bac6b5;
sos_loop[0].somModel.sram_ptr[4][124]=3;
sos_loop[0].somModel.sram_dat[4][125][0]=96'h262308ed;
sos_loop[0].somModel.sram_ptr[4][125]=3;
sos_loop[0].somModel.sram_dat[4][126][0]=96'h82928ac6;
sos_loop[0].somModel.sram_ptr[4][126]=3;
sos_loop[0].somModel.sram_dat[4][127][0]=96'h1fa962b;
sos_loop[0].somModel.sram_ptr[4][127]=3;
sos_loop[0].somModel.sram_dat[4][128][0]=96'h4530cf55;
sos_loop[0].somModel.sram_ptr[4][128]=3;
sos_loop[0].somModel.sram_dat[4][129][0]=96'hb7031fdc;
sos_loop[0].somModel.sram_ptr[4][129]=3;
sos_loop[0].somModel.sram_dat[4][130][0]=96'h3f72ee54;
sos_loop[0].somModel.sram_ptr[4][130]=3;
sos_loop[0].somModel.sram_dat[4][131][0]=96'h4aef92a8;
sos_loop[0].somModel.sram_ptr[4][131]=3;
sos_loop[0].somModel.sram_dat[4][132][0]=96'h7dfb9e62;
sos_loop[0].somModel.sram_ptr[4][132]=3;
sos_loop[0].somModel.sram_dat[4][133][0]=96'hfd4d55c0;
sos_loop[0].somModel.sram_ptr[4][133]=3;
sos_loop[0].somModel.sram_dat[4][134][0]=96'hdf11a902;
sos_loop[0].somModel.sram_ptr[4][134]=3;
sos_loop[0].somModel.sram_dat[4][135][0]=96'ha994cec8;
sos_loop[0].somModel.sram_ptr[4][135]=3;
sos_loop[0].somModel.sram_dat[4][136][0]=96'h8b112348;
sos_loop[0].somModel.sram_ptr[4][136]=3;
sos_loop[0].somModel.sram_dat[4][137][0]=96'hc5b510b9;
sos_loop[0].somModel.sram_ptr[4][137]=3;
sos_loop[0].somModel.sram_dat[4][138][0]=96'h11d4a9aa;
sos_loop[0].somModel.sram_ptr[4][138]=3;
sos_loop[0].somModel.sram_dat[4][139][0]=96'h654037d5;
sos_loop[0].somModel.sram_ptr[4][139]=3;
sos_loop[0].somModel.sram_dat[4][140][0]=96'hb69b89dc;
sos_loop[0].somModel.sram_ptr[4][140]=3;
sos_loop[0].somModel.sram_dat[4][141][0]=96'hd8ece25f;
sos_loop[0].somModel.sram_ptr[4][141]=3;
sos_loop[0].somModel.sram_dat[4][142][0]=96'hef864456;
sos_loop[0].somModel.sram_ptr[4][142]=3;
sos_loop[0].somModel.sram_dat[4][143][0]=96'h7b94efcc;
sos_loop[0].somModel.sram_ptr[4][143]=3;
sos_loop[0].somModel.sram_dat[4][144][0]=96'h5f914f66;
sos_loop[0].somModel.sram_ptr[4][144]=3;
sos_loop[0].somModel.sram_dat[4][145][0]=96'h30cd16e7;
sos_loop[0].somModel.sram_ptr[4][145]=3;
sos_loop[0].somModel.sram_dat[4][146][0]=96'h6e43f380;
sos_loop[0].somModel.sram_ptr[4][146]=3;
sos_loop[0].somModel.sram_dat[4][147][0]=96'haa9b6cac;
sos_loop[0].somModel.sram_ptr[4][147]=3;
sos_loop[0].somModel.sram_dat[4][148][0]=96'hcf4b728d;
sos_loop[0].somModel.sram_ptr[4][148]=3;
sos_loop[0].somModel.sram_dat[4][149][0]=96'h76fbb46a;
sos_loop[0].somModel.sram_ptr[4][149]=3;
sos_loop[0].somModel.sram_dat[4][150][0]=96'h60d90ae;
sos_loop[0].somModel.sram_ptr[4][150]=3;
sos_loop[0].somModel.sram_dat[4][151][0]=96'hcd54a04b;
sos_loop[0].somModel.sram_ptr[4][151]=3;
sos_loop[0].somModel.sram_dat[4][152][0]=96'hcfe265ce;
sos_loop[0].somModel.sram_ptr[4][152]=3;
sos_loop[0].somModel.sram_dat[4][153][0]=96'hf0077206;
sos_loop[0].somModel.sram_ptr[4][153]=3;
sos_loop[0].somModel.sram_dat[4][154][0]=96'h3dd0f100;
sos_loop[0].somModel.sram_ptr[4][154]=3;
sos_loop[0].somModel.sram_dat[4][155][0]=96'hfe370614;
sos_loop[0].somModel.sram_ptr[4][155]=3;
sos_loop[0].somModel.sram_dat[4][156][0]=96'h86391376;
sos_loop[0].somModel.sram_ptr[4][156]=3;
sos_loop[0].somModel.sram_dat[4][157][0]=96'h241d8645;
sos_loop[0].somModel.sram_ptr[4][157]=3;
sos_loop[0].somModel.sram_dat[4][158][0]=96'he054378d;
sos_loop[0].somModel.sram_ptr[4][158]=3;
sos_loop[0].somModel.sram_dat[4][159][0]=96'h584787de;
sos_loop[0].somModel.sram_ptr[4][159]=3;
sos_loop[0].somModel.sram_dat[4][160][0]=96'hc1d8a74;
sos_loop[0].somModel.sram_ptr[4][160]=3;
sos_loop[0].somModel.sram_dat[4][161][0]=96'h8552542f;
sos_loop[0].somModel.sram_ptr[4][161]=3;
sos_loop[0].somModel.sram_dat[4][162][0]=96'h6c061d4c;
sos_loop[0].somModel.sram_ptr[4][162]=3;
sos_loop[0].somModel.sram_dat[4][163][0]=96'h82c410f7;
sos_loop[0].somModel.sram_ptr[4][163]=3;
sos_loop[0].somModel.sram_dat[4][164][0]=96'h1b55f2a5;
sos_loop[0].somModel.sram_ptr[4][164]=3;
sos_loop[0].somModel.sram_dat[4][165][0]=96'h19821382;
sos_loop[0].somModel.sram_ptr[4][165]=3;
sos_loop[0].somModel.sram_dat[4][166][0]=96'hfc383767;
sos_loop[0].somModel.sram_ptr[4][166]=3;
sos_loop[0].somModel.sram_dat[4][167][0]=96'h261dc3a4;
sos_loop[0].somModel.sram_ptr[4][167]=3;
sos_loop[0].somModel.sram_dat[4][168][0]=96'h66ecf2c0;
sos_loop[0].somModel.sram_ptr[4][168]=3;
sos_loop[0].somModel.sram_dat[4][169][0]=96'h52965345;
sos_loop[0].somModel.sram_ptr[4][169]=3;
sos_loop[0].somModel.sram_dat[4][170][0]=96'h33c3d5ba;
sos_loop[0].somModel.sram_ptr[4][170]=3;
sos_loop[0].somModel.sram_dat[4][171][0]=96'h3debd5fc;
sos_loop[0].somModel.sram_ptr[4][171]=3;
sos_loop[0].somModel.sram_dat[4][172][0]=96'h30b16b83;
sos_loop[0].somModel.sram_ptr[4][172]=3;
sos_loop[0].somModel.sram_dat[4][173][0]=96'h9c363d21;
sos_loop[0].somModel.sram_ptr[4][173]=3;
sos_loop[0].somModel.sram_dat[4][174][0]=96'h61a9a8d5;
sos_loop[0].somModel.sram_ptr[4][174]=3;
sos_loop[0].somModel.sram_dat[4][175][0]=96'h7c6464e6;
sos_loop[0].somModel.sram_ptr[4][175]=3;
sos_loop[0].somModel.sram_dat[4][176][0]=96'h122eb0;
sos_loop[0].somModel.sram_ptr[4][176]=3;
sos_loop[0].somModel.sram_dat[4][177][0]=96'h564d3063;
sos_loop[0].somModel.sram_ptr[4][177]=3;
sos_loop[0].somModel.sram_dat[4][178][0]=96'h92ace320;
sos_loop[0].somModel.sram_ptr[4][178]=3;
sos_loop[0].somModel.sram_dat[4][179][0]=96'hd45a4476;
sos_loop[0].somModel.sram_ptr[4][179]=3;
sos_loop[0].somModel.sram_dat[4][180][0]=96'h82700c14;
sos_loop[0].somModel.sram_ptr[4][180]=3;
sos_loop[0].somModel.sram_dat[4][181][0]=96'h51c1fec6;
sos_loop[0].somModel.sram_ptr[4][181]=3;
sos_loop[0].somModel.sram_dat[4][182][0]=96'hbe3dfa7b;
sos_loop[0].somModel.sram_ptr[4][182]=3;
sos_loop[0].somModel.sram_dat[4][183][0]=96'h17e20095;
sos_loop[0].somModel.sram_ptr[4][183]=3;
sos_loop[0].somModel.sram_dat[4][184][0]=96'hd182ec77;
sos_loop[0].somModel.sram_ptr[4][184]=3;
sos_loop[0].somModel.sram_dat[4][185][0]=96'h1917b9b3;
sos_loop[0].somModel.sram_ptr[4][185]=3;
sos_loop[0].somModel.sram_dat[4][186][0]=96'h69a64bf6;
sos_loop[0].somModel.sram_ptr[4][186]=3;
sos_loop[0].somModel.sram_dat[4][187][0]=96'hc48d51a9;
sos_loop[0].somModel.sram_ptr[4][187]=3;
sos_loop[0].somModel.sram_dat[4][188][0]=96'h5a3898ac;
sos_loop[0].somModel.sram_ptr[4][188]=3;
sos_loop[0].somModel.sram_dat[4][189][0]=96'hab1e93a4;
sos_loop[0].somModel.sram_ptr[4][189]=3;
sos_loop[0].somModel.sram_dat[4][190][0]=96'hff34d4ee;
sos_loop[0].somModel.sram_ptr[4][190]=3;
sos_loop[0].somModel.sram_dat[4][191][0]=96'hd7ec1785;
sos_loop[0].somModel.sram_ptr[4][191]=3;
sos_loop[0].somModel.sram_dat[4][192][0]=96'hf631838c;
sos_loop[0].somModel.sram_ptr[4][192]=3;
sos_loop[0].somModel.sram_dat[4][193][0]=96'h70b5c77e;
sos_loop[0].somModel.sram_ptr[4][193]=3;
sos_loop[0].somModel.sram_dat[4][194][0]=96'hf75cba4e;
sos_loop[0].somModel.sram_ptr[4][194]=3;
sos_loop[0].somModel.sram_dat[4][195][0]=96'haa1de942;
sos_loop[0].somModel.sram_ptr[4][195]=3;
sos_loop[0].somModel.sram_dat[4][196][0]=96'h81a5c739;
sos_loop[0].somModel.sram_ptr[4][196]=3;
sos_loop[0].somModel.sram_dat[4][197][0]=96'h99781523;
sos_loop[0].somModel.sram_ptr[4][197]=3;
sos_loop[0].somModel.sram_dat[4][198][0]=96'h728f2c47;
sos_loop[0].somModel.sram_ptr[4][198]=3;
sos_loop[0].somModel.sram_dat[4][199][0]=96'hcaf6348c;
sos_loop[0].somModel.sram_ptr[4][199]=3;
sos_loop[0].somModel.sram_dat[4][200][0]=96'hea9c6e6a;
sos_loop[0].somModel.sram_ptr[4][200]=3;
sos_loop[0].somModel.sram_dat[4][201][0]=96'h29f7a8b6;
sos_loop[0].somModel.sram_ptr[4][201]=3;
sos_loop[0].somModel.sram_dat[4][202][0]=96'hb2b48afc;
sos_loop[0].somModel.sram_ptr[4][202]=3;
sos_loop[0].somModel.sram_dat[4][203][0]=96'h7ce2de;
sos_loop[0].somModel.sram_ptr[4][203]=3;
sos_loop[0].somModel.sram_dat[4][204][0]=96'he9399dcc;
sos_loop[0].somModel.sram_ptr[4][204]=3;
sos_loop[0].somModel.sram_dat[4][205][0]=96'h42d77ee9;
sos_loop[0].somModel.sram_ptr[4][205]=3;
sos_loop[0].somModel.sram_dat[4][206][0]=96'h3fbab7ac;
sos_loop[0].somModel.sram_ptr[4][206]=3;
sos_loop[0].somModel.sram_dat[4][207][0]=96'hd2447ab1;
sos_loop[0].somModel.sram_ptr[4][207]=3;
sos_loop[0].somModel.sram_dat[4][208][0]=96'h1153bd56;
sos_loop[0].somModel.sram_ptr[4][208]=3;
sos_loop[0].somModel.sram_dat[4][209][0]=96'h903d6fbe;
sos_loop[0].somModel.sram_ptr[4][209]=3;
sos_loop[0].somModel.sram_dat[4][210][0]=96'h57510c1;
sos_loop[0].somModel.sram_ptr[4][210]=3;
sos_loop[0].somModel.sram_dat[4][211][0]=96'he6ed5c85;
sos_loop[0].somModel.sram_ptr[4][211]=3;
sos_loop[0].somModel.sram_dat[4][212][0]=96'h311ca0be;
sos_loop[0].somModel.sram_ptr[4][212]=3;
sos_loop[0].somModel.sram_dat[4][213][0]=96'hf7280a93;
sos_loop[0].somModel.sram_ptr[4][213]=3;
sos_loop[0].somModel.sram_dat[4][214][0]=96'h2e6b5b5c;
sos_loop[0].somModel.sram_ptr[4][214]=3;
sos_loop[0].somModel.sram_dat[4][215][0]=96'h46919b60;
sos_loop[0].somModel.sram_ptr[4][215]=3;
sos_loop[0].somModel.sram_dat[4][216][0]=96'hc582966e;
sos_loop[0].somModel.sram_ptr[4][216]=3;
sos_loop[0].somModel.sram_dat[4][217][0]=96'h994201b4;
sos_loop[0].somModel.sram_ptr[4][217]=3;
sos_loop[0].somModel.sram_dat[4][218][0]=96'haa59313;
sos_loop[0].somModel.sram_ptr[4][218]=3;
sos_loop[0].somModel.sram_dat[4][219][0]=96'hbf51da19;
sos_loop[0].somModel.sram_ptr[4][219]=3;
sos_loop[0].somModel.sram_dat[4][220][0]=96'h18fa858a;
sos_loop[0].somModel.sram_ptr[4][220]=3;
sos_loop[0].somModel.sram_dat[4][221][0]=96'h9af5b012;
sos_loop[0].somModel.sram_ptr[4][221]=3;
sos_loop[0].somModel.sram_dat[4][222][0]=96'hfe2e0794;
sos_loop[0].somModel.sram_ptr[4][222]=3;
sos_loop[0].somModel.sram_dat[4][223][0]=96'h86f6eff0;
sos_loop[0].somModel.sram_ptr[4][223]=3;
sos_loop[0].somModel.sram_dat[4][224][0]=96'h6db30707;
sos_loop[0].somModel.sram_ptr[4][224]=3;
sos_loop[0].somModel.sram_dat[4][225][0]=96'h27042389;
sos_loop[0].somModel.sram_ptr[4][225]=3;
sos_loop[0].somModel.sram_dat[4][226][0]=96'h18914c;
sos_loop[0].somModel.sram_ptr[4][226]=3;
sos_loop[0].somModel.sram_dat[4][227][0]=96'h1fe68bc6;
sos_loop[0].somModel.sram_ptr[4][227]=3;
sos_loop[0].somModel.sram_dat[4][228][0]=96'ha4cd25e8;
sos_loop[0].somModel.sram_ptr[4][228]=3;
sos_loop[0].somModel.sram_dat[4][229][0]=96'h9dd2002e;
sos_loop[0].somModel.sram_ptr[4][229]=3;
sos_loop[0].somModel.sram_dat[4][230][0]=96'hfc0a0251;
sos_loop[0].somModel.sram_ptr[4][230]=3;
sos_loop[0].somModel.sram_dat[4][231][0]=96'h3c00e18b;
sos_loop[0].somModel.sram_ptr[4][231]=3;
sos_loop[0].somModel.sram_dat[4][232][0]=96'h1805c387;
sos_loop[0].somModel.sram_ptr[4][232]=3;
sos_loop[0].somModel.sram_dat[4][233][0]=96'h4f21587a;
sos_loop[0].somModel.sram_ptr[4][233]=3;
sos_loop[0].somModel.sram_dat[4][234][0]=96'h182f28a4;
sos_loop[0].somModel.sram_ptr[4][234]=3;
sos_loop[0].somModel.sram_dat[4][235][0]=96'hd1f512d2;
sos_loop[0].somModel.sram_ptr[4][235]=3;
sos_loop[0].somModel.sram_dat[4][236][0]=96'hb807c52d;
sos_loop[0].somModel.sram_ptr[4][236]=3;
sos_loop[0].somModel.sram_dat[4][237][0]=96'he29931ca;
sos_loop[0].somModel.sram_ptr[4][237]=3;
sos_loop[0].somModel.sram_dat[4][238][0]=96'hace9bab6;
sos_loop[0].somModel.sram_ptr[4][238]=3;
sos_loop[0].somModel.sram_dat[4][239][0]=96'hf553012f;
sos_loop[0].somModel.sram_ptr[4][239]=3;
sos_loop[0].somModel.sram_dat[4][240][0]=96'he71db873;
sos_loop[0].somModel.sram_ptr[4][240]=3;
sos_loop[0].somModel.sram_dat[4][241][0]=96'hfa51e2d7;
sos_loop[0].somModel.sram_ptr[4][241]=3;
sos_loop[0].somModel.sram_dat[4][242][0]=96'ha2049980;
sos_loop[0].somModel.sram_ptr[4][242]=3;
sos_loop[0].somModel.sram_dat[4][243][0]=96'hdcabc03c;
sos_loop[0].somModel.sram_ptr[4][243]=3;
sos_loop[0].somModel.sram_dat[4][244][0]=96'heaba455;
sos_loop[0].somModel.sram_ptr[4][244]=3;
sos_loop[0].somModel.sram_dat[4][245][0]=96'ha03e1c48;
sos_loop[0].somModel.sram_ptr[4][245]=3;
sos_loop[0].somModel.sram_dat[4][246][0]=96'hbd9737aa;
sos_loop[0].somModel.sram_ptr[4][246]=3;
sos_loop[0].somModel.sram_dat[4][247][0]=96'h8d5ce6fa;
sos_loop[0].somModel.sram_ptr[4][247]=3;
sos_loop[0].somModel.sram_dat[4][248][0]=96'ha332a6c7;
sos_loop[0].somModel.sram_ptr[4][248]=3;
sos_loop[0].somModel.sram_dat[4][249][0]=96'hd2d22924;
sos_loop[0].somModel.sram_ptr[4][249]=3;
sos_loop[0].somModel.sram_dat[4][250][0]=96'hdb0b6f34;
sos_loop[0].somModel.sram_ptr[4][250]=3;
sos_loop[0].somModel.sram_dat[4][251][0]=96'h205831d3;
sos_loop[0].somModel.sram_ptr[4][251]=3;
sos_loop[0].somModel.sram_dat[4][252][0]=96'h3423f5ae;
sos_loop[0].somModel.sram_ptr[4][252]=3;
sos_loop[0].somModel.sram_dat[4][253][0]=96'hf69a827f;
sos_loop[0].somModel.sram_ptr[4][253]=3;
sos_loop[0].somModel.sram_dat[4][254][0]=96'hd96cf06f;
sos_loop[0].somModel.sram_ptr[4][254]=3;
sos_loop[0].somModel.sram_dat[4][255][0]=96'hab53b800;
sos_loop[0].somModel.sram_ptr[4][255]=3;
sos_loop[0].somModel.sram_dat[4][256][0]=96'h23b65e4f;
sos_loop[0].somModel.sram_ptr[4][256]=3;
sos_loop[0].somModel.sram_dat[4][257][0]=96'h93aeabfb;
sos_loop[0].somModel.sram_ptr[4][257]=3;
sos_loop[0].somModel.sram_dat[4][258][0]=96'hd6166a86;
sos_loop[0].somModel.sram_ptr[4][258]=3;
sos_loop[0].somModel.sram_dat[4][259][0]=96'h14acd40b;
sos_loop[0].somModel.sram_ptr[4][259]=3;
sos_loop[0].somModel.sram_dat[4][260][0]=96'h70c7ab10;
sos_loop[0].somModel.sram_ptr[4][260]=3;
sos_loop[0].somModel.sram_dat[4][261][0]=96'h85c0749b;
sos_loop[0].somModel.sram_ptr[4][261]=3;
sos_loop[0].somModel.sram_dat[4][262][0]=96'h40e49bc4;
sos_loop[0].somModel.sram_ptr[4][262]=3;
sos_loop[0].somModel.sram_dat[4][263][0]=96'hd33d79e6;
sos_loop[0].somModel.sram_ptr[4][263]=3;
sos_loop[0].somModel.sram_dat[4][264][0]=96'h69bcc50f;
sos_loop[0].somModel.sram_ptr[4][264]=3;
sos_loop[0].somModel.sram_dat[4][265][0]=96'h102d9dfb;
sos_loop[0].somModel.sram_ptr[4][265]=3;
sos_loop[0].somModel.sram_dat[4][266][0]=96'hd9113f9f;
sos_loop[0].somModel.sram_ptr[4][266]=3;
sos_loop[0].somModel.sram_dat[4][267][0]=96'h47b3eb80;
sos_loop[0].somModel.sram_ptr[4][267]=3;
sos_loop[0].somModel.sram_dat[4][268][0]=96'heebaf9d5;
sos_loop[0].somModel.sram_ptr[4][268]=3;
sos_loop[0].somModel.sram_dat[4][269][0]=96'hebf5e752;
sos_loop[0].somModel.sram_ptr[4][269]=3;
sos_loop[0].somModel.sram_dat[4][270][0]=96'hc857f0a1;
sos_loop[0].somModel.sram_ptr[4][270]=3;
sos_loop[0].somModel.sram_dat[4][271][0]=96'h79cedbd6;
sos_loop[0].somModel.sram_ptr[4][271]=3;
sos_loop[0].somModel.sram_dat[4][272][0]=96'h719f8337;
sos_loop[0].somModel.sram_ptr[4][272]=3;
sos_loop[0].somModel.sram_dat[4][273][0]=96'h4932ef53;
sos_loop[0].somModel.sram_ptr[4][273]=3;
sos_loop[0].somModel.sram_dat[4][274][0]=96'h79ea4387;
sos_loop[0].somModel.sram_ptr[4][274]=3;
sos_loop[0].somModel.sram_dat[4][275][0]=96'h74a43cf4;
sos_loop[0].somModel.sram_ptr[4][275]=3;
sos_loop[0].somModel.sram_dat[4][276][0]=96'h4fae7a9c;
sos_loop[0].somModel.sram_ptr[4][276]=3;
sos_loop[0].somModel.sram_dat[4][277][0]=96'h117ccf94;
sos_loop[0].somModel.sram_ptr[4][277]=3;
sos_loop[0].somModel.sram_dat[4][278][0]=96'h2009284c;
sos_loop[0].somModel.sram_ptr[4][278]=3;
sos_loop[0].somModel.sram_dat[4][279][0]=96'hfd97e863;
sos_loop[0].somModel.sram_ptr[4][279]=3;
sos_loop[0].somModel.sram_dat[4][280][0]=96'hb4be0194;
sos_loop[0].somModel.sram_ptr[4][280]=3;
sos_loop[0].somModel.sram_dat[4][281][0]=96'h379a4aab;
sos_loop[0].somModel.sram_ptr[4][281]=3;
sos_loop[0].somModel.sram_dat[4][282][0]=96'h19c749de;
sos_loop[0].somModel.sram_ptr[4][282]=3;
sos_loop[0].somModel.sram_dat[4][283][0]=96'h409fb84d;
sos_loop[0].somModel.sram_ptr[4][283]=3;
sos_loop[0].somModel.sram_dat[4][284][0]=96'h3f53200b;
sos_loop[0].somModel.sram_ptr[4][284]=3;
sos_loop[0].somModel.sram_dat[4][285][0]=96'hf7160cc5;
sos_loop[0].somModel.sram_ptr[4][285]=3;
sos_loop[0].somModel.sram_dat[4][286][0]=96'hf8145fad;
sos_loop[0].somModel.sram_ptr[4][286]=3;
sos_loop[0].somModel.sram_dat[4][287][0]=96'hd19b7ecd;
sos_loop[0].somModel.sram_ptr[4][287]=3;
sos_loop[0].somModel.sram_dat[4][288][0]=96'hbb9956a;
sos_loop[0].somModel.sram_ptr[4][288]=3;
sos_loop[0].somModel.sram_dat[4][289][0]=96'hbfc2e567;
sos_loop[0].somModel.sram_ptr[4][289]=3;
sos_loop[0].somModel.sram_dat[4][290][0]=96'hefe2da10;
sos_loop[0].somModel.sram_ptr[4][290]=3;
sos_loop[0].somModel.sram_dat[4][291][0]=96'h8359e399;
sos_loop[0].somModel.sram_ptr[4][291]=3;
sos_loop[0].somModel.sram_dat[4][292][0]=96'h8352ddc5;
sos_loop[0].somModel.sram_ptr[4][292]=3;
sos_loop[0].somModel.sram_dat[4][293][0]=96'h9a537628;
sos_loop[0].somModel.sram_ptr[4][293]=3;
sos_loop[0].somModel.sram_dat[4][294][0]=96'he7259ec5;
sos_loop[0].somModel.sram_ptr[4][294]=3;
sos_loop[0].somModel.sram_dat[4][295][0]=96'ha2aa7d6d;
sos_loop[0].somModel.sram_ptr[4][295]=3;
sos_loop[0].somModel.sram_dat[4][296][0]=96'h562cb1c9;
sos_loop[0].somModel.sram_ptr[4][296]=3;
sos_loop[0].somModel.sram_dat[4][297][0]=96'hf3c4a8d4;
sos_loop[0].somModel.sram_ptr[4][297]=3;
sos_loop[0].somModel.sram_dat[4][298][0]=96'h92ab903f;
sos_loop[0].somModel.sram_ptr[4][298]=3;
sos_loop[0].somModel.sram_dat[4][299][0]=96'h55f5e147;
sos_loop[0].somModel.sram_ptr[4][299]=3;
sos_loop[0].somModel.sram_dat[4][300][0]=96'h7a4d1421;
sos_loop[0].somModel.sram_ptr[4][300]=3;
sos_loop[0].somModel.sram_dat[4][301][0]=96'h7295d548;
sos_loop[0].somModel.sram_ptr[4][301]=3;
sos_loop[0].somModel.sram_dat[4][302][0]=96'h4e27af39;
sos_loop[0].somModel.sram_ptr[4][302]=3;
sos_loop[0].somModel.sram_dat[4][303][0]=96'h3cc0f13c;
sos_loop[0].somModel.sram_ptr[4][303]=3;
sos_loop[0].somModel.sram_dat[4][304][0]=96'h80598983;
sos_loop[0].somModel.sram_ptr[4][304]=3;
sos_loop[0].somModel.sram_dat[4][305][0]=96'h3879539;
sos_loop[0].somModel.sram_ptr[4][305]=3;
sos_loop[0].somModel.sram_dat[4][306][0]=96'hc189aa13;
sos_loop[0].somModel.sram_ptr[4][306]=3;
sos_loop[0].somModel.sram_dat[4][307][0]=96'hc9a30d74;
sos_loop[0].somModel.sram_ptr[4][307]=3;
sos_loop[0].somModel.sram_dat[4][308][0]=96'ha560670f;
sos_loop[0].somModel.sram_ptr[4][308]=3;
sos_loop[0].somModel.sram_dat[4][309][0]=96'h7565e7f0;
sos_loop[0].somModel.sram_ptr[4][309]=3;
sos_loop[0].somModel.sram_dat[4][310][0]=96'h629f25ce;
sos_loop[0].somModel.sram_ptr[4][310]=3;
sos_loop[0].somModel.sram_dat[4][311][0]=96'h55a2a3e;
sos_loop[0].somModel.sram_ptr[4][311]=3;
sos_loop[0].somModel.sram_dat[4][312][0]=96'hb0a85a06;
sos_loop[0].somModel.sram_ptr[4][312]=3;
sos_loop[0].somModel.sram_dat[4][313][0]=96'heeefdd01;
sos_loop[0].somModel.sram_ptr[4][313]=3;
sos_loop[0].somModel.sram_dat[4][314][0]=96'h227ae3eb;
sos_loop[0].somModel.sram_ptr[4][314]=3;
sos_loop[0].somModel.sram_dat[4][315][0]=96'h2bbb2043;
sos_loop[0].somModel.sram_ptr[4][315]=3;
sos_loop[0].somModel.sram_dat[4][316][0]=96'h7c6161ba;
sos_loop[0].somModel.sram_ptr[4][316]=3;
sos_loop[0].somModel.sram_dat[4][317][0]=96'h66da02b6;
sos_loop[0].somModel.sram_ptr[4][317]=3;
sos_loop[0].somModel.sram_dat[4][318][0]=96'h2d6e83ce;
sos_loop[0].somModel.sram_ptr[4][318]=3;
sos_loop[0].somModel.sram_dat[4][319][0]=96'h5e0ed5fd;
sos_loop[0].somModel.sram_ptr[4][319]=3;
sos_loop[0].somModel.sram_dat[4][320][0]=96'h4e41522e;
sos_loop[0].somModel.sram_ptr[4][320]=3;
sos_loop[0].somModel.sram_dat[4][321][0]=96'hd651b46b;
sos_loop[0].somModel.sram_ptr[4][321]=3;
sos_loop[0].somModel.sram_dat[4][322][0]=96'h62d1130b;
sos_loop[0].somModel.sram_ptr[4][322]=3;
sos_loop[0].somModel.sram_dat[4][323][0]=96'hd35fc028;
sos_loop[0].somModel.sram_ptr[4][323]=3;
sos_loop[0].somModel.sram_dat[4][324][0]=96'h5f77f850;
sos_loop[0].somModel.sram_ptr[4][324]=3;
sos_loop[0].somModel.sram_dat[4][325][0]=96'hf6d659f8;
sos_loop[0].somModel.sram_ptr[4][325]=3;
sos_loop[0].somModel.sram_dat[4][326][0]=96'h55963f23;
sos_loop[0].somModel.sram_ptr[4][326]=3;
sos_loop[0].somModel.sram_dat[4][327][0]=96'hd4b3416;
sos_loop[0].somModel.sram_ptr[4][327]=3;
sos_loop[0].somModel.sram_dat[4][328][0]=96'h115c174c;
sos_loop[0].somModel.sram_ptr[4][328]=3;
sos_loop[0].somModel.sram_dat[4][329][0]=96'hc120820c;
sos_loop[0].somModel.sram_ptr[4][329]=3;
sos_loop[0].somModel.sram_dat[4][330][0]=96'hf26eb020;
sos_loop[0].somModel.sram_ptr[4][330]=3;
sos_loop[0].somModel.sram_dat[4][331][0]=96'h13329e53;
sos_loop[0].somModel.sram_ptr[4][331]=3;
sos_loop[0].somModel.sram_dat[4][332][0]=96'h5b10314d;
sos_loop[0].somModel.sram_ptr[4][332]=3;
sos_loop[0].somModel.sram_dat[4][333][0]=96'h1e060ea5;
sos_loop[0].somModel.sram_ptr[4][333]=3;
sos_loop[0].somModel.sram_dat[4][334][0]=96'hff71e09f;
sos_loop[0].somModel.sram_ptr[4][334]=3;
sos_loop[0].somModel.sram_dat[4][335][0]=96'h1f6052ef;
sos_loop[0].somModel.sram_ptr[4][335]=3;
sos_loop[0].somModel.sram_dat[4][336][0]=96'he74d7298;
sos_loop[0].somModel.sram_ptr[4][336]=3;
sos_loop[0].somModel.sram_dat[4][337][0]=96'h6bc68533;
sos_loop[0].somModel.sram_ptr[4][337]=3;
sos_loop[0].somModel.sram_dat[4][338][0]=96'hac2f4971;
sos_loop[0].somModel.sram_ptr[4][338]=3;
sos_loop[0].somModel.sram_dat[4][339][0]=96'he09c405c;
sos_loop[0].somModel.sram_ptr[4][339]=3;
sos_loop[0].somModel.sram_dat[4][340][0]=96'hbbcf571;
sos_loop[0].somModel.sram_ptr[4][340]=3;
sos_loop[0].somModel.sram_dat[4][341][0]=96'h9cb2baa9;
sos_loop[0].somModel.sram_ptr[4][341]=3;
sos_loop[0].somModel.sram_dat[4][342][0]=96'hf9c5b3ea;
sos_loop[0].somModel.sram_ptr[4][342]=3;
sos_loop[0].somModel.sram_dat[4][343][0]=96'hf650f3be;
sos_loop[0].somModel.sram_ptr[4][343]=3;
sos_loop[0].somModel.sram_dat[4][344][0]=96'hd22e73ae;
sos_loop[0].somModel.sram_ptr[4][344]=3;
sos_loop[0].somModel.sram_dat[4][345][0]=96'hd96940ac;
sos_loop[0].somModel.sram_ptr[4][345]=3;
sos_loop[0].somModel.sram_dat[4][346][0]=96'h70cd97c2;
sos_loop[0].somModel.sram_ptr[4][346]=3;
sos_loop[0].somModel.sram_dat[4][347][0]=96'h313273e5;
sos_loop[0].somModel.sram_ptr[4][347]=3;
sos_loop[0].somModel.sram_dat[4][348][0]=96'he79d22d3;
sos_loop[0].somModel.sram_ptr[4][348]=3;
sos_loop[0].somModel.sram_dat[4][349][0]=96'h4542cf7e;
sos_loop[0].somModel.sram_ptr[4][349]=3;
sos_loop[0].somModel.sram_dat[4][350][0]=96'h86391c8b;
sos_loop[0].somModel.sram_ptr[4][350]=3;
sos_loop[0].somModel.sram_dat[4][351][0]=96'h3d91212e;
sos_loop[0].somModel.sram_ptr[4][351]=3;
sos_loop[0].somModel.sram_dat[4][352][0]=96'hc9c85bde;
sos_loop[0].somModel.sram_ptr[4][352]=3;
sos_loop[0].somModel.sram_dat[4][353][0]=96'hc7acf9d9;
sos_loop[0].somModel.sram_ptr[4][353]=3;
sos_loop[0].somModel.sram_dat[4][354][0]=96'hca0ddcf5;
sos_loop[0].somModel.sram_ptr[4][354]=3;
sos_loop[0].somModel.sram_dat[4][355][0]=96'hd10700da;
sos_loop[0].somModel.sram_ptr[4][355]=3;
sos_loop[0].somModel.sram_dat[4][356][0]=96'h3d5daf6b;
sos_loop[0].somModel.sram_ptr[4][356]=3;
sos_loop[0].somModel.sram_dat[4][357][0]=96'h16276984;
sos_loop[0].somModel.sram_ptr[4][357]=3;
sos_loop[0].somModel.sram_dat[4][358][0]=96'h1267258a;
sos_loop[0].somModel.sram_ptr[4][358]=3;
sos_loop[0].somModel.sram_dat[4][359][0]=96'ha7935c99;
sos_loop[0].somModel.sram_ptr[4][359]=3;
sos_loop[0].somModel.sram_dat[4][360][0]=96'h40d7269d;
sos_loop[0].somModel.sram_ptr[4][360]=3;
sos_loop[0].somModel.sram_dat[4][361][0]=96'h3b7070ca;
sos_loop[0].somModel.sram_ptr[4][361]=3;
sos_loop[0].somModel.sram_dat[4][362][0]=96'ha265004e;
sos_loop[0].somModel.sram_ptr[4][362]=3;
sos_loop[0].somModel.sram_dat[4][363][0]=96'h5aa3264;
sos_loop[0].somModel.sram_ptr[4][363]=3;
sos_loop[0].somModel.sram_dat[4][364][0]=96'hfc21ce68;
sos_loop[0].somModel.sram_ptr[4][364]=3;
sos_loop[0].somModel.sram_dat[4][365][0]=96'hee6756c9;
sos_loop[0].somModel.sram_ptr[4][365]=3;
sos_loop[0].somModel.sram_dat[4][366][0]=96'h250a4770;
sos_loop[0].somModel.sram_ptr[4][366]=3;
sos_loop[0].somModel.sram_dat[4][367][0]=96'hbb4715f1;
sos_loop[0].somModel.sram_ptr[4][367]=3;
sos_loop[0].somModel.sram_dat[4][368][0]=96'h257f8471;
sos_loop[0].somModel.sram_ptr[4][368]=3;
sos_loop[0].somModel.sram_dat[4][369][0]=96'h181e4032;
sos_loop[0].somModel.sram_ptr[4][369]=3;
sos_loop[0].somModel.sram_dat[4][370][0]=96'heba8beed;
sos_loop[0].somModel.sram_ptr[4][370]=3;
sos_loop[0].somModel.sram_dat[4][371][0]=96'h550cbdfd;
sos_loop[0].somModel.sram_ptr[4][371]=3;
sos_loop[0].somModel.sram_dat[4][372][0]=96'h312fd6e0;
sos_loop[0].somModel.sram_ptr[4][372]=3;
sos_loop[0].somModel.sram_dat[4][373][0]=96'h51244eaf;
sos_loop[0].somModel.sram_ptr[4][373]=3;
sos_loop[0].somModel.sram_dat[4][374][0]=96'h33bdf527;
sos_loop[0].somModel.sram_ptr[4][374]=3;
sos_loop[0].somModel.sram_dat[4][375][0]=96'hd14622c5;
sos_loop[0].somModel.sram_ptr[4][375]=3;
sos_loop[0].somModel.sram_dat[4][376][0]=96'hdc47ec5f;
sos_loop[0].somModel.sram_ptr[4][376]=3;
sos_loop[0].somModel.sram_dat[4][377][0]=96'h59ac3723;
sos_loop[0].somModel.sram_ptr[4][377]=3;
sos_loop[0].somModel.sram_dat[4][378][0]=96'hc1e60747;
sos_loop[0].somModel.sram_ptr[4][378]=3;
sos_loop[0].somModel.sram_dat[4][379][0]=96'hf7a199f9;
sos_loop[0].somModel.sram_ptr[4][379]=3;
sos_loop[0].somModel.sram_dat[4][380][0]=96'h5bca9a2b;
sos_loop[0].somModel.sram_ptr[4][380]=3;
sos_loop[0].somModel.sram_dat[4][381][0]=96'hd94adb5f;
sos_loop[0].somModel.sram_ptr[4][381]=3;
sos_loop[0].somModel.sram_dat[4][382][0]=96'h9cc28bec;
sos_loop[0].somModel.sram_ptr[4][382]=3;
sos_loop[0].somModel.sram_dat[4][383][0]=96'hf7e9401f;
sos_loop[0].somModel.sram_ptr[4][383]=3;
sos_loop[0].somModel.sram_dat[4][384][0]=96'hc81e26e4;
sos_loop[0].somModel.sram_ptr[4][384]=3;
sos_loop[0].somModel.sram_dat[4][385][0]=96'h3da918ad;
sos_loop[0].somModel.sram_ptr[4][385]=3;
sos_loop[0].somModel.sram_dat[4][386][0]=96'h53f821b7;
sos_loop[0].somModel.sram_ptr[4][386]=3;
sos_loop[0].somModel.sram_dat[4][387][0]=96'he7e00d8b;
sos_loop[0].somModel.sram_ptr[4][387]=3;
sos_loop[0].somModel.sram_dat[4][388][0]=96'h98e3e8fe;
sos_loop[0].somModel.sram_ptr[4][388]=3;
sos_loop[0].somModel.sram_dat[4][389][0]=96'hd66f9e32;
sos_loop[0].somModel.sram_ptr[4][389]=3;
sos_loop[0].somModel.sram_dat[4][390][0]=96'h8afc2cc8;
sos_loop[0].somModel.sram_ptr[4][390]=3;
sos_loop[0].somModel.sram_dat[4][391][0]=96'hdb57684a;
sos_loop[0].somModel.sram_ptr[4][391]=3;
sos_loop[0].somModel.sram_dat[4][392][0]=96'h7f3dad18;
sos_loop[0].somModel.sram_ptr[4][392]=3;
sos_loop[0].somModel.sram_dat[4][393][0]=96'h4a9968a9;
sos_loop[0].somModel.sram_ptr[4][393]=3;
sos_loop[0].somModel.sram_dat[4][394][0]=96'h42710fa3;
sos_loop[0].somModel.sram_ptr[4][394]=3;
sos_loop[0].somModel.sram_dat[4][395][0]=96'h7efb06db;
sos_loop[0].somModel.sram_ptr[4][395]=3;
sos_loop[0].somModel.sram_dat[4][396][0]=96'h958a9fd8;
sos_loop[0].somModel.sram_ptr[4][396]=3;
sos_loop[0].somModel.sram_dat[4][397][0]=96'h6b82013c;
sos_loop[0].somModel.sram_ptr[4][397]=3;
sos_loop[0].somModel.sram_dat[4][398][0]=96'heb6c6952;
sos_loop[0].somModel.sram_ptr[4][398]=3;
sos_loop[0].somModel.sram_dat[4][399][0]=96'h980df882;
sos_loop[0].somModel.sram_ptr[4][399]=3;
sos_loop[0].somModel.sram_dat[4][400][0]=96'h51a3bacd;
sos_loop[0].somModel.sram_ptr[4][400]=3;
sos_loop[0].somModel.sram_dat[4][401][0]=96'hc846112e;
sos_loop[0].somModel.sram_ptr[4][401]=3;
sos_loop[0].somModel.sram_dat[4][402][0]=96'hfbb38c5d;
sos_loop[0].somModel.sram_ptr[4][402]=3;
sos_loop[0].somModel.sram_dat[4][403][0]=96'he94cf512;
sos_loop[0].somModel.sram_ptr[4][403]=3;
sos_loop[0].somModel.sram_dat[4][404][0]=96'hba51e5ae;
sos_loop[0].somModel.sram_ptr[4][404]=3;
sos_loop[0].somModel.sram_dat[4][405][0]=96'h202827f4;
sos_loop[0].somModel.sram_ptr[4][405]=3;
sos_loop[0].somModel.sram_dat[4][406][0]=96'hf29e4104;
sos_loop[0].somModel.sram_ptr[4][406]=3;
sos_loop[0].somModel.sram_dat[4][407][0]=96'h7644bccf;
sos_loop[0].somModel.sram_ptr[4][407]=3;
sos_loop[0].somModel.sram_dat[4][408][0]=96'hdd35657;
sos_loop[0].somModel.sram_ptr[4][408]=3;
sos_loop[0].somModel.sram_dat[4][409][0]=96'h415386ed;
sos_loop[0].somModel.sram_ptr[4][409]=3;
sos_loop[0].somModel.sram_dat[4][410][0]=96'h3576469;
sos_loop[0].somModel.sram_ptr[4][410]=3;
sos_loop[0].somModel.sram_dat[4][411][0]=96'h1fbc279b;
sos_loop[0].somModel.sram_ptr[4][411]=3;
sos_loop[0].somModel.sram_dat[4][412][0]=96'ha271cab3;
sos_loop[0].somModel.sram_ptr[4][412]=3;
sos_loop[0].somModel.sram_dat[4][413][0]=96'h712d2a8d;
sos_loop[0].somModel.sram_ptr[4][413]=3;
sos_loop[0].somModel.sram_dat[4][414][0]=96'h3fddf6b3;
sos_loop[0].somModel.sram_ptr[4][414]=3;
sos_loop[0].somModel.sram_dat[4][415][0]=96'h2165be7a;
sos_loop[0].somModel.sram_ptr[4][415]=3;
sos_loop[0].somModel.sram_dat[4][416][0]=96'h448d049b;
sos_loop[0].somModel.sram_ptr[4][416]=3;
sos_loop[0].somModel.sram_dat[4][417][0]=96'hfb2d5087;
sos_loop[0].somModel.sram_ptr[4][417]=3;
sos_loop[0].somModel.sram_dat[4][418][0]=96'h1e98ac81;
sos_loop[0].somModel.sram_ptr[4][418]=3;
sos_loop[0].somModel.sram_dat[4][419][0]=96'he671ad3e;
sos_loop[0].somModel.sram_ptr[4][419]=3;
sos_loop[0].somModel.sram_dat[4][420][0]=96'hc5704dd4;
sos_loop[0].somModel.sram_ptr[4][420]=3;
sos_loop[0].somModel.sram_dat[4][421][0]=96'hb0840ac8;
sos_loop[0].somModel.sram_ptr[4][421]=3;
sos_loop[0].somModel.sram_dat[4][422][0]=96'hfa0d4b7c;
sos_loop[0].somModel.sram_ptr[4][422]=3;
sos_loop[0].somModel.sram_dat[4][423][0]=96'hea1183e1;
sos_loop[0].somModel.sram_ptr[4][423]=3;
sos_loop[0].somModel.sram_dat[4][424][0]=96'hb91fade1;
sos_loop[0].somModel.sram_ptr[4][424]=3;
sos_loop[0].somModel.sram_dat[4][425][0]=96'ha11fde54;
sos_loop[0].somModel.sram_ptr[4][425]=3;
sos_loop[0].somModel.sram_dat[4][426][0]=96'h12eff59c;
sos_loop[0].somModel.sram_ptr[4][426]=3;
sos_loop[0].somModel.sram_dat[4][427][0]=96'hdb238c5d;
sos_loop[0].somModel.sram_ptr[4][427]=3;
sos_loop[0].somModel.sram_dat[4][428][0]=96'hc55954a;
sos_loop[0].somModel.sram_ptr[4][428]=3;
sos_loop[0].somModel.sram_dat[4][429][0]=96'h4160f5ee;
sos_loop[0].somModel.sram_ptr[4][429]=3;
sos_loop[0].somModel.sram_dat[4][430][0]=96'hedcbd779;
sos_loop[0].somModel.sram_ptr[4][430]=3;
sos_loop[0].somModel.sram_dat[4][431][0]=96'hf4a82895;
sos_loop[0].somModel.sram_ptr[4][431]=3;
sos_loop[0].somModel.sram_dat[4][432][0]=96'h1604c030;
sos_loop[0].somModel.sram_ptr[4][432]=3;
sos_loop[0].somModel.sram_dat[4][433][0]=96'hc0a439bf;
sos_loop[0].somModel.sram_ptr[4][433]=3;
sos_loop[0].somModel.sram_dat[4][434][0]=96'h2a955aec;
sos_loop[0].somModel.sram_ptr[4][434]=3;
sos_loop[0].somModel.sram_dat[4][435][0]=96'h2c902099;
sos_loop[0].somModel.sram_ptr[4][435]=3;
sos_loop[0].somModel.sram_dat[4][436][0]=96'h217c7717;
sos_loop[0].somModel.sram_ptr[4][436]=3;
sos_loop[0].somModel.sram_dat[4][437][0]=96'h7c0ea408;
sos_loop[0].somModel.sram_ptr[4][437]=3;
sos_loop[0].somModel.sram_dat[4][438][0]=96'h4d0afc5c;
sos_loop[0].somModel.sram_ptr[4][438]=3;
sos_loop[0].somModel.sram_dat[4][439][0]=96'hb8cd0eab;
sos_loop[0].somModel.sram_ptr[4][439]=3;
sos_loop[0].somModel.sram_dat[4][440][0]=96'h739e2b20;
sos_loop[0].somModel.sram_ptr[4][440]=3;
sos_loop[0].somModel.sram_dat[4][441][0]=96'h34dbf565;
sos_loop[0].somModel.sram_ptr[4][441]=3;
sos_loop[0].somModel.sram_dat[4][442][0]=96'h66f2d912;
sos_loop[0].somModel.sram_ptr[4][442]=3;
sos_loop[0].somModel.sram_dat[4][443][0]=96'hb7295d4e;
sos_loop[0].somModel.sram_ptr[4][443]=3;
sos_loop[0].somModel.sram_dat[4][444][0]=96'h316d5676;
sos_loop[0].somModel.sram_ptr[4][444]=3;
sos_loop[0].somModel.sram_dat[4][445][0]=96'h69aa0de2;
sos_loop[0].somModel.sram_ptr[4][445]=3;
sos_loop[0].somModel.sram_dat[4][446][0]=96'h7110b17d;
sos_loop[0].somModel.sram_ptr[4][446]=3;
sos_loop[0].somModel.sram_dat[4][447][0]=96'h93b4e0f7;
sos_loop[0].somModel.sram_ptr[4][447]=3;
sos_loop[0].somModel.sram_dat[4][448][0]=96'h4dc5b038;
sos_loop[0].somModel.sram_ptr[4][448]=3;
sos_loop[0].somModel.sram_dat[4][449][0]=96'hb9e03453;
sos_loop[0].somModel.sram_ptr[4][449]=3;
sos_loop[0].somModel.sram_dat[4][450][0]=96'hf831c057;
sos_loop[0].somModel.sram_ptr[4][450]=3;
sos_loop[0].somModel.sram_dat[4][451][0]=96'h3834ff31;
sos_loop[0].somModel.sram_ptr[4][451]=3;
sos_loop[0].somModel.sram_dat[4][452][0]=96'hbcbc82bf;
sos_loop[0].somModel.sram_ptr[4][452]=3;
sos_loop[0].somModel.sram_dat[4][453][0]=96'h4c1bec8b;
sos_loop[0].somModel.sram_ptr[4][453]=3;
sos_loop[0].somModel.sram_dat[4][454][0]=96'h209ec751;
sos_loop[0].somModel.sram_ptr[4][454]=3;
sos_loop[0].somModel.sram_dat[4][455][0]=96'h4de18e05;
sos_loop[0].somModel.sram_ptr[4][455]=3;
sos_loop[0].somModel.sram_dat[4][456][0]=96'h4f7ba449;
sos_loop[0].somModel.sram_ptr[4][456]=3;
sos_loop[0].somModel.sram_dat[4][457][0]=96'h6036359;
sos_loop[0].somModel.sram_ptr[4][457]=3;
sos_loop[0].somModel.sram_dat[4][458][0]=96'h712983c2;
sos_loop[0].somModel.sram_ptr[4][458]=3;
sos_loop[0].somModel.sram_dat[4][459][0]=96'h20770d60;
sos_loop[0].somModel.sram_ptr[4][459]=3;
sos_loop[0].somModel.sram_dat[4][460][0]=96'hf63206a4;
sos_loop[0].somModel.sram_ptr[4][460]=3;
sos_loop[0].somModel.sram_dat[4][461][0]=96'h72a80a04;
sos_loop[0].somModel.sram_ptr[4][461]=3;
sos_loop[0].somModel.sram_dat[4][462][0]=96'hd8d85182;
sos_loop[0].somModel.sram_ptr[4][462]=3;
sos_loop[0].somModel.sram_dat[4][463][0]=96'h965e1956;
sos_loop[0].somModel.sram_ptr[4][463]=3;
sos_loop[0].somModel.sram_dat[4][464][0]=96'h71bce5d1;
sos_loop[0].somModel.sram_ptr[4][464]=3;
sos_loop[0].somModel.sram_dat[4][465][0]=96'h1acccf4d;
sos_loop[0].somModel.sram_ptr[4][465]=3;
sos_loop[0].somModel.sram_dat[4][466][0]=96'hbe3c6600;
sos_loop[0].somModel.sram_ptr[4][466]=3;
sos_loop[0].somModel.sram_dat[4][467][0]=96'hf6b42162;
sos_loop[0].somModel.sram_ptr[4][467]=3;
sos_loop[0].somModel.sram_dat[4][468][0]=96'h1ebef7e4;
sos_loop[0].somModel.sram_ptr[4][468]=3;
sos_loop[0].somModel.sram_dat[4][469][0]=96'h449b815e;
sos_loop[0].somModel.sram_ptr[4][469]=3;
sos_loop[0].somModel.sram_dat[4][470][0]=96'hf700305c;
sos_loop[0].somModel.sram_ptr[4][470]=3;
sos_loop[0].somModel.sram_dat[4][471][0]=96'h71d16c63;
sos_loop[0].somModel.sram_ptr[4][471]=3;
sos_loop[0].somModel.sram_dat[4][472][0]=96'haf7769e2;
sos_loop[0].somModel.sram_ptr[4][472]=3;
sos_loop[0].somModel.sram_dat[4][473][0]=96'h9238595d;
sos_loop[0].somModel.sram_ptr[4][473]=3;
sos_loop[0].somModel.sram_dat[4][474][0]=96'h87abb692;
sos_loop[0].somModel.sram_ptr[4][474]=3;
sos_loop[0].somModel.sram_dat[4][475][0]=96'h9f619149;
sos_loop[0].somModel.sram_ptr[4][475]=3;
sos_loop[0].somModel.sram_dat[4][476][0]=96'h1c452d06;
sos_loop[0].somModel.sram_ptr[4][476]=3;
sos_loop[0].somModel.sram_dat[4][477][0]=96'h47627aba;
sos_loop[0].somModel.sram_ptr[4][477]=3;
sos_loop[0].somModel.sram_dat[4][478][0]=96'h751c717c;
sos_loop[0].somModel.sram_ptr[4][478]=3;
sos_loop[0].somModel.sram_dat[4][479][0]=96'hca65525a;
sos_loop[0].somModel.sram_ptr[4][479]=3;
sos_loop[0].somModel.sram_dat[4][480][0]=96'hb8645166;
sos_loop[0].somModel.sram_ptr[4][480]=3;
sos_loop[0].somModel.sram_dat[4][481][0]=96'ha9a978fb;
sos_loop[0].somModel.sram_ptr[4][481]=3;
sos_loop[0].somModel.sram_dat[4][482][0]=96'h4f00fbb0;
sos_loop[0].somModel.sram_ptr[4][482]=3;
sos_loop[0].somModel.sram_dat[4][483][0]=96'hdc1e87e7;
sos_loop[0].somModel.sram_ptr[4][483]=3;
sos_loop[0].somModel.sram_dat[4][484][0]=96'h6b81d355;
sos_loop[0].somModel.sram_ptr[4][484]=3;
sos_loop[0].somModel.sram_dat[4][485][0]=96'h3e7fe58b;
sos_loop[0].somModel.sram_ptr[4][485]=3;
sos_loop[0].somModel.sram_dat[4][486][0]=96'hf3f20799;
sos_loop[0].somModel.sram_ptr[4][486]=3;
sos_loop[0].somModel.sram_dat[4][487][0]=96'hc30e1c35;
sos_loop[0].somModel.sram_ptr[4][487]=3;
sos_loop[0].somModel.sram_dat[4][488][0]=96'hda9ad8a1;
sos_loop[0].somModel.sram_ptr[4][488]=3;
sos_loop[0].somModel.sram_dat[4][489][0]=96'hfa5f7769;
sos_loop[0].somModel.sram_ptr[4][489]=3;
sos_loop[0].somModel.sram_dat[4][490][0]=96'hb1447c06;
sos_loop[0].somModel.sram_ptr[4][490]=3;
sos_loop[0].somModel.sram_dat[4][491][0]=96'hf95a7eb1;
sos_loop[0].somModel.sram_ptr[4][491]=3;
sos_loop[0].somModel.sram_dat[4][492][0]=96'h9391d306;
sos_loop[0].somModel.sram_ptr[4][492]=3;
sos_loop[0].somModel.sram_dat[4][493][0]=96'h699e2b00;
sos_loop[0].somModel.sram_ptr[4][493]=3;
sos_loop[0].somModel.sram_dat[4][494][0]=96'h891868ba;
sos_loop[0].somModel.sram_ptr[4][494]=3;
sos_loop[0].somModel.sram_dat[4][495][0]=96'ha2b05c48;
sos_loop[0].somModel.sram_ptr[4][495]=3;
sos_loop[0].somModel.sram_dat[4][496][0]=96'haac8ca5a;
sos_loop[0].somModel.sram_ptr[4][496]=3;
sos_loop[0].somModel.sram_dat[4][497][0]=96'h5f8471bd;
sos_loop[0].somModel.sram_ptr[4][497]=3;
sos_loop[0].somModel.sram_dat[4][498][0]=96'hd0610bc;
sos_loop[0].somModel.sram_ptr[4][498]=3;
sos_loop[0].somModel.sram_dat[4][499][0]=96'h18206fc9;
sos_loop[0].somModel.sram_ptr[4][499]=3;
sos_loop[0].somModel.sram_dat[4][500][0]=96'hac2f36d;
sos_loop[0].somModel.sram_ptr[4][500]=3;
sos_loop[0].somModel.sram_dat[4][501][0]=96'h2e748e8;
sos_loop[0].somModel.sram_ptr[4][501]=3;
sos_loop[0].somModel.sram_dat[4][502][0]=96'hf11fb9e2;
sos_loop[0].somModel.sram_ptr[4][502]=3;
sos_loop[0].somModel.sram_dat[4][503][0]=96'h5b9ea50a;
sos_loop[0].somModel.sram_ptr[4][503]=3;
sos_loop[0].somModel.sram_dat[4][504][0]=96'hf227c657;
sos_loop[0].somModel.sram_ptr[4][504]=3;
sos_loop[0].somModel.sram_dat[4][505][0]=96'h3515ab3b;
sos_loop[0].somModel.sram_ptr[4][505]=3;
sos_loop[0].somModel.sram_dat[4][506][0]=96'h15503f8d;
sos_loop[0].somModel.sram_ptr[4][506]=3;
sos_loop[0].somModel.sram_dat[4][507][0]=96'h76cc4124;
sos_loop[0].somModel.sram_ptr[4][507]=3;
sos_loop[0].somModel.sram_dat[4][508][0]=96'hd4bdec61;
sos_loop[0].somModel.sram_ptr[4][508]=3;
sos_loop[0].somModel.sram_dat[4][509][0]=96'hd2bd71db;
sos_loop[0].somModel.sram_ptr[4][509]=3;
sos_loop[0].somModel.sram_dat[4][510][0]=96'he0a2b56f;
sos_loop[0].somModel.sram_ptr[4][510]=3;
sos_loop[0].somModel.sram_dat[4][511][0]=96'he34d64c6;
sos_loop[0].somModel.sram_ptr[4][511]=3;
sos_loop[0].somModel.sram_dat[4][512][0]=96'hc735ad48;
sos_loop[0].somModel.sram_ptr[4][512]=3;
sos_loop[0].somModel.sram_dat[4][513][0]=96'h7035214f;
sos_loop[0].somModel.sram_ptr[4][513]=3;
sos_loop[0].somModel.sram_dat[4][514][0]=96'hd2ff291a;
sos_loop[0].somModel.sram_ptr[4][514]=3;
sos_loop[0].somModel.sram_dat[4][515][0]=96'h49b6cb18;
sos_loop[0].somModel.sram_ptr[4][515]=3;
sos_loop[0].somModel.sram_dat[4][516][0]=96'hc6cd4467;
sos_loop[0].somModel.sram_ptr[4][516]=3;
sos_loop[0].somModel.sram_dat[4][517][0]=96'he90fe281;
sos_loop[0].somModel.sram_ptr[4][517]=3;
sos_loop[0].somModel.sram_dat[4][518][0]=96'hba02a11d;
sos_loop[0].somModel.sram_ptr[4][518]=3;
sos_loop[0].somModel.sram_dat[4][519][0]=96'h253c7a3;
sos_loop[0].somModel.sram_ptr[4][519]=3;
sos_loop[0].somModel.sram_dat[4][520][0]=96'h412bb30c;
sos_loop[0].somModel.sram_ptr[4][520]=3;
sos_loop[0].somModel.sram_dat[4][521][0]=96'h8d12dd56;
sos_loop[0].somModel.sram_ptr[4][521]=3;
sos_loop[0].somModel.sram_dat[4][522][0]=96'h6fe0c5a1;
sos_loop[0].somModel.sram_ptr[4][522]=3;
sos_loop[0].somModel.sram_dat[4][523][0]=96'ha33b35e9;
sos_loop[0].somModel.sram_ptr[4][523]=3;
sos_loop[0].somModel.sram_dat[4][524][0]=96'h723a31b7;
sos_loop[0].somModel.sram_ptr[4][524]=3;
sos_loop[0].somModel.sram_dat[4][525][0]=96'h5a350d96;
sos_loop[0].somModel.sram_ptr[4][525]=3;
sos_loop[0].somModel.sram_dat[4][526][0]=96'h4006207;
sos_loop[0].somModel.sram_ptr[4][526]=3;
sos_loop[0].somModel.sram_dat[4][527][0]=96'hc702e976;
sos_loop[0].somModel.sram_ptr[4][527]=3;
sos_loop[0].somModel.sram_dat[4][528][0]=96'hb6010e92;
sos_loop[0].somModel.sram_ptr[4][528]=3;
sos_loop[0].somModel.sram_dat[4][529][0]=96'h4c85212;
sos_loop[0].somModel.sram_ptr[4][529]=3;
sos_loop[0].somModel.sram_dat[4][530][0]=96'h40044411;
sos_loop[0].somModel.sram_ptr[4][530]=3;
sos_loop[0].somModel.sram_dat[4][531][0]=96'ha8fb5d85;
sos_loop[0].somModel.sram_ptr[4][531]=3;
sos_loop[0].somModel.sram_dat[4][532][0]=96'h4d9741f6;
sos_loop[0].somModel.sram_ptr[4][532]=3;
sos_loop[0].somModel.sram_dat[4][533][0]=96'hd3afd823;
sos_loop[0].somModel.sram_ptr[4][533]=3;
sos_loop[0].somModel.sram_dat[4][534][0]=96'hfdd6ea42;
sos_loop[0].somModel.sram_ptr[4][534]=3;
sos_loop[0].somModel.sram_dat[4][535][0]=96'hb42b3094;
sos_loop[0].somModel.sram_ptr[4][535]=3;
sos_loop[0].somModel.sram_dat[4][536][0]=96'h2b35ac93;
sos_loop[0].somModel.sram_ptr[4][536]=3;
sos_loop[0].somModel.sram_dat[4][537][0]=96'h1de14302;
sos_loop[0].somModel.sram_ptr[4][537]=3;
sos_loop[0].somModel.sram_dat[4][538][0]=96'h197646ab;
sos_loop[0].somModel.sram_ptr[4][538]=3;
sos_loop[0].somModel.sram_dat[4][539][0]=96'hc205d69;
sos_loop[0].somModel.sram_ptr[4][539]=3;
sos_loop[0].somModel.sram_dat[4][540][0]=96'h8947a1d6;
sos_loop[0].somModel.sram_ptr[4][540]=3;
sos_loop[0].somModel.sram_dat[4][541][0]=96'h6890668;
sos_loop[0].somModel.sram_ptr[4][541]=3;
sos_loop[0].somModel.sram_dat[4][542][0]=96'h8bdb4cbe;
sos_loop[0].somModel.sram_ptr[4][542]=3;
sos_loop[0].somModel.sram_dat[4][543][0]=96'h1969b688;
sos_loop[0].somModel.sram_ptr[4][543]=3;
sos_loop[0].somModel.sram_dat[4][544][0]=96'h10e2ee9c;
sos_loop[0].somModel.sram_ptr[4][544]=3;
sos_loop[0].somModel.sram_dat[4][545][0]=96'ha7e49978;
sos_loop[0].somModel.sram_ptr[4][545]=3;
sos_loop[0].somModel.sram_dat[4][546][0]=96'h860c996f;
sos_loop[0].somModel.sram_ptr[4][546]=3;
sos_loop[0].somModel.sram_dat[4][547][0]=96'hbe168c0d;
sos_loop[0].somModel.sram_ptr[4][547]=3;
sos_loop[0].somModel.sram_dat[4][548][0]=96'hf9cf89b1;
sos_loop[0].somModel.sram_ptr[4][548]=3;
sos_loop[0].somModel.sram_dat[4][549][0]=96'h81261f85;
sos_loop[0].somModel.sram_ptr[4][549]=3;
sos_loop[0].somModel.sram_dat[4][550][0]=96'he7aaa8fd;
sos_loop[0].somModel.sram_ptr[4][550]=3;
sos_loop[0].somModel.sram_dat[4][551][0]=96'hb0429c43;
sos_loop[0].somModel.sram_ptr[4][551]=3;
sos_loop[0].somModel.sram_dat[4][552][0]=96'h8a4c6218;
sos_loop[0].somModel.sram_ptr[4][552]=3;
sos_loop[0].somModel.sram_dat[4][553][0]=96'h95f19822;
sos_loop[0].somModel.sram_ptr[4][553]=3;
sos_loop[0].somModel.sram_dat[4][554][0]=96'h45858f52;
sos_loop[0].somModel.sram_ptr[4][554]=3;
sos_loop[0].somModel.sram_dat[4][555][0]=96'hd544fa47;
sos_loop[0].somModel.sram_ptr[4][555]=3;
sos_loop[0].somModel.sram_dat[4][556][0]=96'haf1a4005;
sos_loop[0].somModel.sram_ptr[4][556]=3;
sos_loop[0].somModel.sram_dat[4][557][0]=96'he3b732bb;
sos_loop[0].somModel.sram_ptr[4][557]=3;
sos_loop[0].somModel.sram_dat[4][558][0]=96'h6194cbd6;
sos_loop[0].somModel.sram_ptr[4][558]=3;
sos_loop[0].somModel.sram_dat[4][559][0]=96'h9d1b6b4b;
sos_loop[0].somModel.sram_ptr[4][559]=3;
sos_loop[0].somModel.sram_dat[4][560][0]=96'h2ff0666f;
sos_loop[0].somModel.sram_ptr[4][560]=3;
sos_loop[0].somModel.sram_dat[4][561][0]=96'h6913bb5f;
sos_loop[0].somModel.sram_ptr[4][561]=3;
sos_loop[0].somModel.sram_dat[4][562][0]=96'h4925a9b2;
sos_loop[0].somModel.sram_ptr[4][562]=3;
sos_loop[0].somModel.sram_dat[4][563][0]=96'hcbf76125;
sos_loop[0].somModel.sram_ptr[4][563]=3;
sos_loop[0].somModel.sram_dat[4][564][0]=96'h80f0a6a3;
sos_loop[0].somModel.sram_ptr[4][564]=3;
sos_loop[0].somModel.sram_dat[4][565][0]=96'h1249cd1d;
sos_loop[0].somModel.sram_ptr[4][565]=3;
sos_loop[0].somModel.sram_dat[4][566][0]=96'hbc0a568e;
sos_loop[0].somModel.sram_ptr[4][566]=3;
sos_loop[0].somModel.sram_dat[4][567][0]=96'h688f87cd;
sos_loop[0].somModel.sram_ptr[4][567]=3;
sos_loop[0].somModel.sram_dat[4][568][0]=96'h2960aaef;
sos_loop[0].somModel.sram_ptr[4][568]=3;
sos_loop[0].somModel.sram_dat[4][569][0]=96'h5085236f;
sos_loop[0].somModel.sram_ptr[4][569]=3;
sos_loop[0].somModel.sram_dat[4][570][0]=96'hef5d2004;
sos_loop[0].somModel.sram_ptr[4][570]=3;
sos_loop[0].somModel.sram_dat[4][571][0]=96'h25b2c4aa;
sos_loop[0].somModel.sram_ptr[4][571]=3;
sos_loop[0].somModel.sram_dat[4][572][0]=96'hb972ba2f;
sos_loop[0].somModel.sram_ptr[4][572]=3;
sos_loop[0].somModel.sram_dat[4][573][0]=96'hfb315574;
sos_loop[0].somModel.sram_ptr[4][573]=3;
sos_loop[0].somModel.sram_dat[4][574][0]=96'h4874d5e7;
sos_loop[0].somModel.sram_ptr[4][574]=3;
sos_loop[0].somModel.sram_dat[4][575][0]=96'h8dfdecc3;
sos_loop[0].somModel.sram_ptr[4][575]=3;
sos_loop[0].somModel.sram_dat[4][576][0]=96'hcce699ec;
sos_loop[0].somModel.sram_ptr[4][576]=3;
sos_loop[0].somModel.sram_dat[4][577][0]=96'h785b1a49;
sos_loop[0].somModel.sram_ptr[4][577]=3;
sos_loop[0].somModel.sram_dat[4][578][0]=96'hebe00791;
sos_loop[0].somModel.sram_ptr[4][578]=3;
sos_loop[0].somModel.sram_dat[4][579][0]=96'hc3beb879;
sos_loop[0].somModel.sram_ptr[4][579]=3;
sos_loop[0].somModel.sram_dat[4][580][0]=96'he4c31860;
sos_loop[0].somModel.sram_ptr[4][580]=3;
sos_loop[0].somModel.sram_dat[4][581][0]=96'hd6fbba7;
sos_loop[0].somModel.sram_ptr[4][581]=3;
sos_loop[0].somModel.sram_dat[4][582][0]=96'hf165457d;
sos_loop[0].somModel.sram_ptr[4][582]=3;
sos_loop[0].somModel.sram_dat[4][583][0]=96'h3805f41d;
sos_loop[0].somModel.sram_ptr[4][583]=3;
sos_loop[0].somModel.sram_dat[4][584][0]=96'h58045c79;
sos_loop[0].somModel.sram_ptr[4][584]=3;
sos_loop[0].somModel.sram_dat[4][585][0]=96'hb77beed9;
sos_loop[0].somModel.sram_ptr[4][585]=3;
sos_loop[0].somModel.sram_dat[4][586][0]=96'h364e16c5;
sos_loop[0].somModel.sram_ptr[4][586]=3;
sos_loop[0].somModel.sram_dat[4][587][0]=96'h379023ab;
sos_loop[0].somModel.sram_ptr[4][587]=3;
sos_loop[0].somModel.sram_dat[4][588][0]=96'h1f3f2a95;
sos_loop[0].somModel.sram_ptr[4][588]=3;
sos_loop[0].somModel.sram_dat[4][589][0]=96'h6317bf23;
sos_loop[0].somModel.sram_ptr[4][589]=3;
sos_loop[0].somModel.sram_dat[4][590][0]=96'h75d392b5;
sos_loop[0].somModel.sram_ptr[4][590]=3;
sos_loop[0].somModel.sram_dat[4][591][0]=96'hd7f4bb13;
sos_loop[0].somModel.sram_ptr[4][591]=3;
sos_loop[0].somModel.sram_dat[4][592][0]=96'hbdf1b95a;
sos_loop[0].somModel.sram_ptr[4][592]=3;
sos_loop[0].somModel.sram_dat[4][593][0]=96'hff3fdc47;
sos_loop[0].somModel.sram_ptr[4][593]=3;
sos_loop[0].somModel.sram_dat[4][594][0]=96'hfe817339;
sos_loop[0].somModel.sram_ptr[4][594]=3;
sos_loop[0].somModel.sram_dat[4][595][0]=96'hb670bd6a;
sos_loop[0].somModel.sram_ptr[4][595]=3;
sos_loop[0].somModel.sram_dat[4][596][0]=96'h80fb1afb;
sos_loop[0].somModel.sram_ptr[4][596]=3;
sos_loop[0].somModel.sram_dat[4][597][0]=96'h7e488471;
sos_loop[0].somModel.sram_ptr[4][597]=3;
sos_loop[0].somModel.sram_dat[4][598][0]=96'h180ab825;
sos_loop[0].somModel.sram_ptr[4][598]=3;
sos_loop[0].somModel.sram_dat[4][599][0]=96'h432afc9f;
sos_loop[0].somModel.sram_ptr[4][599]=3;
sos_loop[0].somModel.sram_dat[4][600][0]=96'he23107c;
sos_loop[0].somModel.sram_ptr[4][600]=3;
sos_loop[0].somModel.sram_dat[4][601][0]=96'h266062f1;
sos_loop[0].somModel.sram_ptr[4][601]=3;
sos_loop[0].somModel.sram_dat[4][602][0]=96'h2ff8a855;
sos_loop[0].somModel.sram_ptr[4][602]=3;
sos_loop[0].somModel.sram_dat[4][603][0]=96'h1ba59a2e;
sos_loop[0].somModel.sram_ptr[4][603]=3;
sos_loop[0].somModel.sram_dat[4][604][0]=96'h3a0d39c7;
sos_loop[0].somModel.sram_ptr[4][604]=3;
sos_loop[0].somModel.sram_dat[4][605][0]=96'h98c7b823;
sos_loop[0].somModel.sram_ptr[4][605]=3;
sos_loop[0].somModel.sram_dat[4][606][0]=96'h5462a053;
sos_loop[0].somModel.sram_ptr[4][606]=3;
sos_loop[0].somModel.sram_dat[4][607][0]=96'hced324b2;
sos_loop[0].somModel.sram_ptr[4][607]=3;
sos_loop[0].somModel.sram_dat[4][608][0]=96'h7808026c;
sos_loop[0].somModel.sram_ptr[4][608]=3;
sos_loop[0].somModel.sram_dat[4][609][0]=96'h76544554;
sos_loop[0].somModel.sram_ptr[4][609]=3;
sos_loop[0].somModel.sram_dat[4][610][0]=96'h587748f1;
sos_loop[0].somModel.sram_ptr[4][610]=3;
sos_loop[0].somModel.sram_dat[4][611][0]=96'hf759b497;
sos_loop[0].somModel.sram_ptr[4][611]=3;
sos_loop[0].somModel.sram_dat[4][612][0]=96'h49dd7a37;
sos_loop[0].somModel.sram_ptr[4][612]=3;
sos_loop[0].somModel.sram_dat[4][613][0]=96'hb16968b0;
sos_loop[0].somModel.sram_ptr[4][613]=3;
sos_loop[0].somModel.sram_dat[4][614][0]=96'h80c27aff;
sos_loop[0].somModel.sram_ptr[4][614]=3;
sos_loop[0].somModel.sram_dat[4][615][0]=96'hd5249c05;
sos_loop[0].somModel.sram_ptr[4][615]=3;
sos_loop[0].somModel.sram_dat[4][616][0]=96'h9b3bb04a;
sos_loop[0].somModel.sram_ptr[4][616]=3;
sos_loop[0].somModel.sram_dat[4][617][0]=96'hc4f06715;
sos_loop[0].somModel.sram_ptr[4][617]=3;
sos_loop[0].somModel.sram_dat[4][618][0]=96'h60e58984;
sos_loop[0].somModel.sram_ptr[4][618]=3;
sos_loop[0].somModel.sram_dat[4][619][0]=96'ha69c4dec;
sos_loop[0].somModel.sram_ptr[4][619]=3;
sos_loop[0].somModel.sram_dat[4][620][0]=96'h9996b95e;
sos_loop[0].somModel.sram_ptr[4][620]=3;
sos_loop[0].somModel.sram_dat[4][621][0]=96'hb3533b00;
sos_loop[0].somModel.sram_ptr[4][621]=3;
sos_loop[0].somModel.sram_dat[4][622][0]=96'h6034dd18;
sos_loop[0].somModel.sram_ptr[4][622]=3;
sos_loop[0].somModel.sram_dat[4][623][0]=96'h74e86cc8;
sos_loop[0].somModel.sram_ptr[4][623]=3;
sos_loop[0].somModel.sram_dat[4][624][0]=96'ha06c8f64;
sos_loop[0].somModel.sram_ptr[4][624]=3;
sos_loop[0].somModel.sram_dat[4][625][0]=96'h3f2bc9a0;
sos_loop[0].somModel.sram_ptr[4][625]=3;
sos_loop[0].somModel.sram_dat[4][626][0]=96'hf81585e9;
sos_loop[0].somModel.sram_ptr[4][626]=3;
sos_loop[0].somModel.sram_dat[4][627][0]=96'h97515402;
sos_loop[0].somModel.sram_ptr[4][627]=3;
sos_loop[0].somModel.sram_dat[4][628][0]=96'h2a07f05;
sos_loop[0].somModel.sram_ptr[4][628]=3;
sos_loop[0].somModel.sram_dat[4][629][0]=96'h2bc32216;
sos_loop[0].somModel.sram_ptr[4][629]=3;
sos_loop[0].somModel.sram_dat[4][630][0]=96'h909c5b0d;
sos_loop[0].somModel.sram_ptr[4][630]=3;
sos_loop[0].somModel.sram_dat[4][631][0]=96'he5dcf0e6;
sos_loop[0].somModel.sram_ptr[4][631]=3;
sos_loop[0].somModel.sram_dat[4][632][0]=96'h965ce467;
sos_loop[0].somModel.sram_ptr[4][632]=3;
sos_loop[0].somModel.sram_dat[4][633][0]=96'h2fe7f356;
sos_loop[0].somModel.sram_ptr[4][633]=3;
sos_loop[0].somModel.sram_dat[4][634][0]=96'h30d25e12;
sos_loop[0].somModel.sram_ptr[4][634]=3;
sos_loop[0].somModel.sram_dat[4][635][0]=96'h4bb8ac18;
sos_loop[0].somModel.sram_ptr[4][635]=3;
sos_loop[0].somModel.sram_dat[4][636][0]=96'h44f4a58a;
sos_loop[0].somModel.sram_ptr[4][636]=3;
sos_loop[0].somModel.sram_dat[4][637][0]=96'hf501287;
sos_loop[0].somModel.sram_ptr[4][637]=3;
sos_loop[0].somModel.sram_dat[4][638][0]=96'h7eaf6d4f;
sos_loop[0].somModel.sram_ptr[4][638]=3;
sos_loop[0].somModel.sram_dat[4][639][0]=96'hd82212f1;
sos_loop[0].somModel.sram_ptr[4][639]=3;
sos_loop[0].somModel.sram_dat[4][640][0]=96'hec1625ea;
sos_loop[0].somModel.sram_ptr[4][640]=3;
sos_loop[0].somModel.sram_dat[4][641][0]=96'h74cae5e1;
sos_loop[0].somModel.sram_ptr[4][641]=3;
sos_loop[0].somModel.sram_dat[4][642][0]=96'h1fe03adc;
sos_loop[0].somModel.sram_ptr[4][642]=3;
sos_loop[0].somModel.sram_dat[4][643][0]=96'he0ce0e82;
sos_loop[0].somModel.sram_ptr[4][643]=3;
sos_loop[0].somModel.sram_dat[4][644][0]=96'h5f82b623;
sos_loop[0].somModel.sram_ptr[4][644]=3;
sos_loop[0].somModel.sram_dat[4][645][0]=96'h7e2be26;
sos_loop[0].somModel.sram_ptr[4][645]=3;
sos_loop[0].somModel.sram_dat[4][646][0]=96'hb4c4d344;
sos_loop[0].somModel.sram_ptr[4][646]=3;
sos_loop[0].somModel.sram_dat[4][647][0]=96'h2ecd929;
sos_loop[0].somModel.sram_ptr[4][647]=3;
sos_loop[0].somModel.sram_dat[4][648][0]=96'hc583cf7b;
sos_loop[0].somModel.sram_ptr[4][648]=3;
sos_loop[0].somModel.sram_dat[4][649][0]=96'hf4373181;
sos_loop[0].somModel.sram_ptr[4][649]=3;
sos_loop[0].somModel.sram_dat[4][650][0]=96'hc69ba9fb;
sos_loop[0].somModel.sram_ptr[4][650]=3;
sos_loop[0].somModel.sram_dat[4][651][0]=96'h8b43e12f;
sos_loop[0].somModel.sram_ptr[4][651]=3;
sos_loop[0].somModel.sram_dat[4][652][0]=96'h1a7a8797;
sos_loop[0].somModel.sram_ptr[4][652]=3;
sos_loop[0].somModel.sram_dat[4][653][0]=96'h6dcbaa62;
sos_loop[0].somModel.sram_ptr[4][653]=3;
sos_loop[0].somModel.sram_dat[4][654][0]=96'h46285e0;
sos_loop[0].somModel.sram_ptr[4][654]=3;
sos_loop[0].somModel.sram_dat[4][655][0]=96'hc9e05443;
sos_loop[0].somModel.sram_ptr[4][655]=3;
sos_loop[0].somModel.sram_dat[4][656][0]=96'h7f136176;
sos_loop[0].somModel.sram_ptr[4][656]=3;
sos_loop[0].somModel.sram_dat[4][657][0]=96'ha9a396f;
sos_loop[0].somModel.sram_ptr[4][657]=3;
sos_loop[0].somModel.sram_dat[4][658][0]=96'hd535e00d;
sos_loop[0].somModel.sram_ptr[4][658]=3;
sos_loop[0].somModel.sram_dat[4][659][0]=96'h76394b0c;
sos_loop[0].somModel.sram_ptr[4][659]=3;
sos_loop[0].somModel.sram_dat[4][660][0]=96'ha330561;
sos_loop[0].somModel.sram_ptr[4][660]=3;
sos_loop[0].somModel.sram_dat[4][661][0]=96'h43b01a49;
sos_loop[0].somModel.sram_ptr[4][661]=3;
sos_loop[0].somModel.sram_dat[4][662][0]=96'hff999355;
sos_loop[0].somModel.sram_ptr[4][662]=3;
sos_loop[0].somModel.sram_dat[4][663][0]=96'ha5eddcfb;
sos_loop[0].somModel.sram_ptr[4][663]=3;
sos_loop[0].somModel.sram_dat[4][664][0]=96'h45f82b33;
sos_loop[0].somModel.sram_ptr[4][664]=3;
sos_loop[0].somModel.sram_dat[4][665][0]=96'h4a4c1e12;
sos_loop[0].somModel.sram_ptr[4][665]=3;
sos_loop[0].somModel.sram_dat[4][666][0]=96'h3b8a6857;
sos_loop[0].somModel.sram_ptr[4][666]=3;
sos_loop[0].somModel.sram_dat[4][667][0]=96'hb1e16a4c;
sos_loop[0].somModel.sram_ptr[4][667]=3;
sos_loop[0].somModel.sram_dat[4][668][0]=96'hfce324ac;
sos_loop[0].somModel.sram_ptr[4][668]=3;
sos_loop[0].somModel.sram_dat[4][669][0]=96'he619bc20;
sos_loop[0].somModel.sram_ptr[4][669]=3;
sos_loop[0].somModel.sram_dat[4][670][0]=96'h2caded6b;
sos_loop[0].somModel.sram_ptr[4][670]=3;
sos_loop[0].somModel.sram_dat[4][671][0]=96'h3b50576b;
sos_loop[0].somModel.sram_ptr[4][671]=3;
sos_loop[0].somModel.sram_dat[4][672][0]=96'h640ef1ce;
sos_loop[0].somModel.sram_ptr[4][672]=3;
sos_loop[0].somModel.sram_dat[4][673][0]=96'hf21564b1;
sos_loop[0].somModel.sram_ptr[4][673]=3;
sos_loop[0].somModel.sram_dat[4][674][0]=96'h25f779da;
sos_loop[0].somModel.sram_ptr[4][674]=3;
sos_loop[0].somModel.sram_dat[4][675][0]=96'h425844e1;
sos_loop[0].somModel.sram_ptr[4][675]=3;
sos_loop[0].somModel.sram_dat[4][676][0]=96'he8c91e81;
sos_loop[0].somModel.sram_ptr[4][676]=3;
sos_loop[0].somModel.sram_dat[4][677][0]=96'h8c9c6fa7;
sos_loop[0].somModel.sram_ptr[4][677]=3;
sos_loop[0].somModel.sram_dat[4][678][0]=96'h79a69237;
sos_loop[0].somModel.sram_ptr[4][678]=3;
sos_loop[0].somModel.sram_dat[4][679][0]=96'h1db22a87;
sos_loop[0].somModel.sram_ptr[4][679]=3;
sos_loop[0].somModel.sram_dat[4][680][0]=96'h243c5486;
sos_loop[0].somModel.sram_ptr[4][680]=3;
sos_loop[0].somModel.sram_dat[4][681][0]=96'h935fc3ce;
sos_loop[0].somModel.sram_ptr[4][681]=3;
sos_loop[0].somModel.sram_dat[4][682][0]=96'h590e4270;
sos_loop[0].somModel.sram_ptr[4][682]=3;
sos_loop[0].somModel.sram_dat[4][683][0]=96'h707e28f6;
sos_loop[0].somModel.sram_ptr[4][683]=3;
sos_loop[0].somModel.sram_dat[4][684][0]=96'hdae57a3d;
sos_loop[0].somModel.sram_ptr[4][684]=3;
sos_loop[0].somModel.sram_dat[4][685][0]=96'hb87638d9;
sos_loop[0].somModel.sram_ptr[4][685]=3;
sos_loop[0].somModel.sram_dat[4][686][0]=96'hd4807ce9;
sos_loop[0].somModel.sram_ptr[4][686]=3;
sos_loop[0].somModel.sram_dat[4][687][0]=96'h8c9c8a90;
sos_loop[0].somModel.sram_ptr[4][687]=3;
sos_loop[0].somModel.sram_dat[4][688][0]=96'h785a9702;
sos_loop[0].somModel.sram_ptr[4][688]=3;
sos_loop[0].somModel.sram_dat[4][689][0]=96'hb1259e5a;
sos_loop[0].somModel.sram_ptr[4][689]=3;
sos_loop[0].somModel.sram_dat[4][690][0]=96'h9cb6c8e9;
sos_loop[0].somModel.sram_ptr[4][690]=3;
sos_loop[0].somModel.sram_dat[4][691][0]=96'h641e0603;
sos_loop[0].somModel.sram_ptr[4][691]=3;
sos_loop[0].somModel.sram_dat[4][692][0]=96'hfa391441;
sos_loop[0].somModel.sram_ptr[4][692]=3;
sos_loop[0].somModel.sram_dat[4][693][0]=96'h2b6458e0;
sos_loop[0].somModel.sram_ptr[4][693]=3;
sos_loop[0].somModel.sram_dat[4][694][0]=96'h268cf6b2;
sos_loop[0].somModel.sram_ptr[4][694]=3;
sos_loop[0].somModel.sram_dat[4][695][0]=96'h7858cb29;
sos_loop[0].somModel.sram_ptr[4][695]=3;
sos_loop[0].somModel.sram_dat[4][696][0]=96'hc0447d97;
sos_loop[0].somModel.sram_ptr[4][696]=3;
sos_loop[0].somModel.sram_dat[4][697][0]=96'habd5331;
sos_loop[0].somModel.sram_ptr[4][697]=3;
sos_loop[0].somModel.sram_dat[4][698][0]=96'h8ccb7b91;
sos_loop[0].somModel.sram_ptr[4][698]=3;
sos_loop[0].somModel.sram_dat[4][699][0]=96'h722790a4;
sos_loop[0].somModel.sram_ptr[4][699]=3;
sos_loop[0].somModel.sram_dat[4][700][0]=96'h1de04b8;
sos_loop[0].somModel.sram_ptr[4][700]=3;
sos_loop[0].somModel.cfg_tbl_sel[4] = 4;
sos_loop[0].somModel.cfg_dat_sel[4] = 3;
sos_loop[0].somModel.cfg_dat_vld[4] = 1;
sos_loop[0].somModel.cfg_miss_ptr[4] = 0;
sos_loop[0].somModel.tcam_data[5][0][0]=80'h00000000000000000000;
sos_loop[0].somModel.tcam_mask[5][0][0]=80'hffffffffffffffffffff;
sos_loop[0].somModel.tcam_data[5][1][0]=80'h00000000c76428a3ac18;
sos_loop[0].somModel.tcam_mask[5][1][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][2][0]=80'h000000006fa2b332a044;
sos_loop[0].somModel.tcam_mask[5][2][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][3][0]=80'h00000000df160ea7e244;
sos_loop[0].somModel.tcam_mask[5][3][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][4][0]=80'h00000000bde8a5158a2b;
sos_loop[0].somModel.tcam_mask[5][4][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][5][0]=80'h000000001c7fcaa5772f;
sos_loop[0].somModel.tcam_mask[5][5][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][6][0]=80'h00000000398bc2065413;
sos_loop[0].somModel.tcam_mask[5][6][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][7][0]=80'h00000000bf26a132d23e;
sos_loop[0].somModel.tcam_mask[5][7][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][8][0]=80'h000000002e5a52ddfb3f;
sos_loop[0].somModel.tcam_mask[5][8][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][9][0]=80'h000000000f9c4f448c4c;
sos_loop[0].somModel.tcam_mask[5][9][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][10][0]=80'h0000000035e4dd182f90;
sos_loop[0].somModel.tcam_mask[5][10][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][11][0]=80'h000000008513d0c50521;
sos_loop[0].somModel.tcam_mask[5][11][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][12][0]=80'h0000000035a66285b62e;
sos_loop[0].somModel.tcam_mask[5][12][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][13][0]=80'h000000004915d9de428f;
sos_loop[0].somModel.tcam_mask[5][13][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][14][0]=80'h000000003eff489073c2;
sos_loop[0].somModel.tcam_mask[5][14][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][15][0]=80'h00000000d00165db49c5;
sos_loop[0].somModel.tcam_mask[5][15][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][16][0]=80'h00000000c6e7d540048a;
sos_loop[0].somModel.tcam_mask[5][16][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][17][0]=80'h000000000d2cf31221e9;
sos_loop[0].somModel.tcam_mask[5][17][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][18][0]=80'h000000009cc2400c08bc;
sos_loop[0].somModel.tcam_mask[5][18][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][19][0]=80'h00000000e84ab68b1a24;
sos_loop[0].somModel.tcam_mask[5][19][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][20][0]=80'h00000000dc9c606e91ae;
sos_loop[0].somModel.tcam_mask[5][20][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][21][0]=80'h000000004b8ee53f7660;
sos_loop[0].somModel.tcam_mask[5][21][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][22][0]=80'h00000000a6dc109cdbbd;
sos_loop[0].somModel.tcam_mask[5][22][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][23][0]=80'h000000002e5acd726cb2;
sos_loop[0].somModel.tcam_mask[5][23][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][24][0]=80'h00000000bb30b2ecd487;
sos_loop[0].somModel.tcam_mask[5][24][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][25][0]=80'h000000009aeec82f8fac;
sos_loop[0].somModel.tcam_mask[5][25][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][26][0]=80'h00000000ab83fe2b985c;
sos_loop[0].somModel.tcam_mask[5][26][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][27][0]=80'h00000000ca3daac02b2f;
sos_loop[0].somModel.tcam_mask[5][27][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][28][0]=80'h000000001a893b2ffa10;
sos_loop[0].somModel.tcam_mask[5][28][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][29][0]=80'h00000000cb1ab883d9ca;
sos_loop[0].somModel.tcam_mask[5][29][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][30][0]=80'h000000006ddb0412e88d;
sos_loop[0].somModel.tcam_mask[5][30][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][31][0]=80'h0000000025d034a677c8;
sos_loop[0].somModel.tcam_mask[5][31][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][32][0]=80'h0000000002ee63ce89af;
sos_loop[0].somModel.tcam_mask[5][32][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[5][33][0]=80'h000000001ab5a710d843;
sos_loop[0].somModel.tcam_mask[5][33][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][34][0]=80'h0000000097e8c062f084;
sos_loop[0].somModel.tcam_mask[5][34][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][35][0]=80'h0000000030a809743d4f;
sos_loop[0].somModel.tcam_mask[5][35][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][36][0]=80'h0000000022420da7f8f4;
sos_loop[0].somModel.tcam_mask[5][36][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][37][0]=80'h00000000afaf284ad3bc;
sos_loop[0].somModel.tcam_mask[5][37][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][38][0]=80'h0000000053bd4f0d7794;
sos_loop[0].somModel.tcam_mask[5][38][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][39][0]=80'h000000005c0d39f2f061;
sos_loop[0].somModel.tcam_mask[5][39][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][40][0]=80'h000000009419a7ce074a;
sos_loop[0].somModel.tcam_mask[5][40][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][41][0]=80'h00000000052d45cc1e4a;
sos_loop[0].somModel.tcam_mask[5][41][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][42][0]=80'h000000009b30665b9971;
sos_loop[0].somModel.tcam_mask[5][42][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][43][0]=80'h0000000020d936f412c1;
sos_loop[0].somModel.tcam_mask[5][43][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][44][0]=80'h000000008b889af41550;
sos_loop[0].somModel.tcam_mask[5][44][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][45][0]=80'h00000000f91ce85e797d;
sos_loop[0].somModel.tcam_mask[5][45][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][46][0]=80'h0000000006e1dbd81191;
sos_loop[0].somModel.tcam_mask[5][46][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][47][0]=80'h00000000345e3c5f1365;
sos_loop[0].somModel.tcam_mask[5][47][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][48][0]=80'h000000008dceefe91dc9;
sos_loop[0].somModel.tcam_mask[5][48][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][49][0]=80'h00000000d47d2191ffed;
sos_loop[0].somModel.tcam_mask[5][49][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][50][0]=80'h000000007d341fbc821b;
sos_loop[0].somModel.tcam_mask[5][50][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][51][0]=80'h000000002e1c5d9ff7d9;
sos_loop[0].somModel.tcam_mask[5][51][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][52][0]=80'h00000000b7c667fd0324;
sos_loop[0].somModel.tcam_mask[5][52][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][53][0]=80'h000000004933bf21a16c;
sos_loop[0].somModel.tcam_mask[5][53][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][54][0]=80'h00000000f9724902347e;
sos_loop[0].somModel.tcam_mask[5][54][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][55][0]=80'h00000000aeb766b220db;
sos_loop[0].somModel.tcam_mask[5][55][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][56][0]=80'h00000000dbbc2a3224ab;
sos_loop[0].somModel.tcam_mask[5][56][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][57][0]=80'h00000000365a679e8085;
sos_loop[0].somModel.tcam_mask[5][57][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][58][0]=80'h00000000eeff7c2b7b33;
sos_loop[0].somModel.tcam_mask[5][58][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][59][0]=80'h0000000045bb6a31bb68;
sos_loop[0].somModel.tcam_mask[5][59][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][60][0]=80'h000000001a81b1c43f91;
sos_loop[0].somModel.tcam_mask[5][60][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][61][0]=80'h000000001de0ad29184a;
sos_loop[0].somModel.tcam_mask[5][61][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][62][0]=80'h000000004eb9229cd415;
sos_loop[0].somModel.tcam_mask[5][62][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][63][0]=80'h0000000075c39cfd15db;
sos_loop[0].somModel.tcam_mask[5][63][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][64][0]=80'h000000000bd7d9ddf726;
sos_loop[0].somModel.tcam_mask[5][64][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][65][0]=80'h00000000788ece7eed43;
sos_loop[0].somModel.tcam_mask[5][65][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][66][0]=80'h00000000689790000fff;
sos_loop[0].somModel.tcam_mask[5][66][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][67][0]=80'h0000000030fca31cf96b;
sos_loop[0].somModel.tcam_mask[5][67][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][68][0]=80'h00000000358975cc2823;
sos_loop[0].somModel.tcam_mask[5][68][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][69][0]=80'h000000006b1cd921c79d;
sos_loop[0].somModel.tcam_mask[5][69][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][70][0]=80'h00000000549a31ff63b7;
sos_loop[0].somModel.tcam_mask[5][70][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][71][0]=80'h00000000310dee607220;
sos_loop[0].somModel.tcam_mask[5][71][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][72][0]=80'h00000000af90fc2fb606;
sos_loop[0].somModel.tcam_mask[5][72][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][73][0]=80'h000000000db655000d3a;
sos_loop[0].somModel.tcam_mask[5][73][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][74][0]=80'h000000008bf35344ab45;
sos_loop[0].somModel.tcam_mask[5][74][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][75][0]=80'h000000002d8a38190b20;
sos_loop[0].somModel.tcam_mask[5][75][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][76][0]=80'h000000000263f7f66582;
sos_loop[0].somModel.tcam_mask[5][76][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[5][77][0]=80'h000000004dfc2ba4768d;
sos_loop[0].somModel.tcam_mask[5][77][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][78][0]=80'h00000000849983bfbe7a;
sos_loop[0].somModel.tcam_mask[5][78][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][79][0]=80'h000000001efcb2f4dd4d;
sos_loop[0].somModel.tcam_mask[5][79][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][80][0]=80'h0000000061e5a9de4569;
sos_loop[0].somModel.tcam_mask[5][80][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][81][0]=80'h00000000770c1c4bd3a5;
sos_loop[0].somModel.tcam_mask[5][81][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][82][0]=80'h00000000500562660aff;
sos_loop[0].somModel.tcam_mask[5][82][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][83][0]=80'h00000000a72a189143e2;
sos_loop[0].somModel.tcam_mask[5][83][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][84][0]=80'h0000000051a64abf0e09;
sos_loop[0].somModel.tcam_mask[5][84][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][85][0]=80'h000000001f5700abe928;
sos_loop[0].somModel.tcam_mask[5][85][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][86][0]=80'h00000000512e72fad6a2;
sos_loop[0].somModel.tcam_mask[5][86][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][87][0]=80'h000000005f3a530396cf;
sos_loop[0].somModel.tcam_mask[5][87][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][88][0]=80'h00000000748487400445;
sos_loop[0].somModel.tcam_mask[5][88][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][89][0]=80'h0000000087719fb3f864;
sos_loop[0].somModel.tcam_mask[5][89][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][90][0]=80'h00000000e88c8f60061d;
sos_loop[0].somModel.tcam_mask[5][90][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][91][0]=80'h000000009f6cc5f93019;
sos_loop[0].somModel.tcam_mask[5][91][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][92][0]=80'h00000000fa9df2c0fa11;
sos_loop[0].somModel.tcam_mask[5][92][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][93][0]=80'h000000003e5de237f4f3;
sos_loop[0].somModel.tcam_mask[5][93][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][94][0]=80'h000000001220e6f8b9fd;
sos_loop[0].somModel.tcam_mask[5][94][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][95][0]=80'h00000000ceb0c2f94c3c;
sos_loop[0].somModel.tcam_mask[5][95][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][96][0]=80'h000000001845b8356ded;
sos_loop[0].somModel.tcam_mask[5][96][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][97][0]=80'h00000000cb7d6f052ed9;
sos_loop[0].somModel.tcam_mask[5][97][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][98][0]=80'h00000000a1d827523dc7;
sos_loop[0].somModel.tcam_mask[5][98][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][99][0]=80'h000000000caf8264a3ea;
sos_loop[0].somModel.tcam_mask[5][99][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][100][0]=80'h0000000038ead3f12916;
sos_loop[0].somModel.tcam_mask[5][100][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][101][0]=80'h0000000013d2ee37c448;
sos_loop[0].somModel.tcam_mask[5][101][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][102][0]=80'h000000003c2fe7d9f34c;
sos_loop[0].somModel.tcam_mask[5][102][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][103][0]=80'h000000003c1db8626079;
sos_loop[0].somModel.tcam_mask[5][103][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][104][0]=80'h00000000865b861ca607;
sos_loop[0].somModel.tcam_mask[5][104][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][105][0]=80'h00000000794600c6d0f4;
sos_loop[0].somModel.tcam_mask[5][105][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][106][0]=80'h00000000e00c57f6e0b3;
sos_loop[0].somModel.tcam_mask[5][106][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][107][0]=80'h00000000e29db65e8903;
sos_loop[0].somModel.tcam_mask[5][107][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][108][0]=80'h000000008e261e6170f3;
sos_loop[0].somModel.tcam_mask[5][108][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][109][0]=80'h0000000066939b10ec73;
sos_loop[0].somModel.tcam_mask[5][109][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][110][0]=80'h0000000070c2e9c3c8eb;
sos_loop[0].somModel.tcam_mask[5][110][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][111][0]=80'h0000000045c66be84cf4;
sos_loop[0].somModel.tcam_mask[5][111][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][112][0]=80'h00000000232cef211d0e;
sos_loop[0].somModel.tcam_mask[5][112][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][113][0]=80'h0000000080542dda5aa2;
sos_loop[0].somModel.tcam_mask[5][113][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][114][0]=80'h00000000474effbc30dd;
sos_loop[0].somModel.tcam_mask[5][114][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][115][0]=80'h00000000e4cebd5c6fa4;
sos_loop[0].somModel.tcam_mask[5][115][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][116][0]=80'h00000000af6a54830375;
sos_loop[0].somModel.tcam_mask[5][116][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][117][0]=80'h000000008ef028be44c1;
sos_loop[0].somModel.tcam_mask[5][117][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][118][0]=80'h000000005fdca8436bf4;
sos_loop[0].somModel.tcam_mask[5][118][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][119][0]=80'h000000006e7e1c15bd08;
sos_loop[0].somModel.tcam_mask[5][119][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][120][0]=80'h00000000134c1f65fd66;
sos_loop[0].somModel.tcam_mask[5][120][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][121][0]=80'h00000000cea87493679f;
sos_loop[0].somModel.tcam_mask[5][121][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][122][0]=80'h00000000ceb7bc309c1a;
sos_loop[0].somModel.tcam_mask[5][122][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][123][0]=80'h0000000061a6f8771878;
sos_loop[0].somModel.tcam_mask[5][123][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][124][0]=80'h00000000cedef6a567fe;
sos_loop[0].somModel.tcam_mask[5][124][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][125][0]=80'h000000002e32a08622cd;
sos_loop[0].somModel.tcam_mask[5][125][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][126][0]=80'h000000005356e16b8fd7;
sos_loop[0].somModel.tcam_mask[5][126][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][127][0]=80'h00000000fd605bd942c3;
sos_loop[0].somModel.tcam_mask[5][127][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][128][0]=80'h0000000000d5f103f449;
sos_loop[0].somModel.tcam_mask[5][128][0]=80'hffffffffff0000000000;
sos_loop[0].somModel.tcam_data[5][129][0]=80'h000000005f57f4362b22;
sos_loop[0].somModel.tcam_mask[5][129][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][130][0]=80'h000000002e67f284f871;
sos_loop[0].somModel.tcam_mask[5][130][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][131][0]=80'h00000000ecd79dcadc01;
sos_loop[0].somModel.tcam_mask[5][131][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][132][0]=80'h00000000e00525c7b0f8;
sos_loop[0].somModel.tcam_mask[5][132][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][133][0]=80'h00000000b3cf483e6c80;
sos_loop[0].somModel.tcam_mask[5][133][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][134][0]=80'h0000000077eb26f31bbe;
sos_loop[0].somModel.tcam_mask[5][134][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][135][0]=80'h000000008b676c49d915;
sos_loop[0].somModel.tcam_mask[5][135][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][136][0]=80'h000000000a2822acbd35;
sos_loop[0].somModel.tcam_mask[5][136][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][137][0]=80'h0000000003a257929df1;
sos_loop[0].somModel.tcam_mask[5][137][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[5][138][0]=80'h00000000e9b0e1c40a18;
sos_loop[0].somModel.tcam_mask[5][138][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][139][0]=80'h000000003f10a0b32f42;
sos_loop[0].somModel.tcam_mask[5][139][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][140][0]=80'h00000000f8a042a8b1d1;
sos_loop[0].somModel.tcam_mask[5][140][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][141][0]=80'h00000000c010041f98fe;
sos_loop[0].somModel.tcam_mask[5][141][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][142][0]=80'h000000006f5155d6bf2a;
sos_loop[0].somModel.tcam_mask[5][142][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][143][0]=80'h000000006174e0aee88e;
sos_loop[0].somModel.tcam_mask[5][143][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][144][0]=80'h00000000d8f296505931;
sos_loop[0].somModel.tcam_mask[5][144][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][145][0]=80'h00000000e512e3c64789;
sos_loop[0].somModel.tcam_mask[5][145][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][146][0]=80'h00000000373e0b9976b9;
sos_loop[0].somModel.tcam_mask[5][146][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][147][0]=80'h0000000003e7dacda18b;
sos_loop[0].somModel.tcam_mask[5][147][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[5][148][0]=80'h000000000964ddbc00a5;
sos_loop[0].somModel.tcam_mask[5][148][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][149][0]=80'h0000000054781b947c65;
sos_loop[0].somModel.tcam_mask[5][149][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][150][0]=80'h000000004e476ae23070;
sos_loop[0].somModel.tcam_mask[5][150][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][151][0]=80'h00000000965a202c5dd1;
sos_loop[0].somModel.tcam_mask[5][151][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][152][0]=80'h000000006eeef25e5a0e;
sos_loop[0].somModel.tcam_mask[5][152][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][153][0]=80'h00000000bd9be825e53c;
sos_loop[0].somModel.tcam_mask[5][153][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][154][0]=80'h000000005a0d2b0e2652;
sos_loop[0].somModel.tcam_mask[5][154][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][155][0]=80'h00000000f02c2960a78f;
sos_loop[0].somModel.tcam_mask[5][155][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][156][0]=80'h0000000043801573ed5c;
sos_loop[0].somModel.tcam_mask[5][156][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][157][0]=80'h0000000034d1a3628645;
sos_loop[0].somModel.tcam_mask[5][157][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][158][0]=80'h00000000476d2c7ebc16;
sos_loop[0].somModel.tcam_mask[5][158][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][159][0]=80'h00000000a17de6c9b9c6;
sos_loop[0].somModel.tcam_mask[5][159][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][160][0]=80'h000000002e3b2da7cb0e;
sos_loop[0].somModel.tcam_mask[5][160][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][161][0]=80'h00000000618fe75b3a00;
sos_loop[0].somModel.tcam_mask[5][161][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][162][0]=80'h000000007868e9b929a2;
sos_loop[0].somModel.tcam_mask[5][162][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][163][0]=80'h00000000cbe5e4137d1a;
sos_loop[0].somModel.tcam_mask[5][163][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][164][0]=80'h000000006771e8c490b5;
sos_loop[0].somModel.tcam_mask[5][164][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][165][0]=80'h000000007be9cc15dbad;
sos_loop[0].somModel.tcam_mask[5][165][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][166][0]=80'h000000008c89b097b14c;
sos_loop[0].somModel.tcam_mask[5][166][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][167][0]=80'h00000000f2124342ae18;
sos_loop[0].somModel.tcam_mask[5][167][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][168][0]=80'h00000000330261ba3670;
sos_loop[0].somModel.tcam_mask[5][168][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][169][0]=80'h0000000042c4edb6d896;
sos_loop[0].somModel.tcam_mask[5][169][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][170][0]=80'h0000000023a570bc32da;
sos_loop[0].somModel.tcam_mask[5][170][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][171][0]=80'h00000000db4f2973fc73;
sos_loop[0].somModel.tcam_mask[5][171][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][172][0]=80'h000000004c40d88318b1;
sos_loop[0].somModel.tcam_mask[5][172][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][173][0]=80'h000000001273739101e3;
sos_loop[0].somModel.tcam_mask[5][173][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][174][0]=80'h000000009c2ebac8770d;
sos_loop[0].somModel.tcam_mask[5][174][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][175][0]=80'h00000000aaeaffde1744;
sos_loop[0].somModel.tcam_mask[5][175][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][176][0]=80'h0000000067b1d0406ac4;
sos_loop[0].somModel.tcam_mask[5][176][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][177][0]=80'h00000000602be7c25423;
sos_loop[0].somModel.tcam_mask[5][177][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][178][0]=80'h000000007bd2374d89da;
sos_loop[0].somModel.tcam_mask[5][178][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][179][0]=80'h00000000484efbf68ee5;
sos_loop[0].somModel.tcam_mask[5][179][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][180][0]=80'h000000008c2970d5df55;
sos_loop[0].somModel.tcam_mask[5][180][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][181][0]=80'h00000000aec65cebfe7b;
sos_loop[0].somModel.tcam_mask[5][181][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][182][0]=80'h0000000094dfc4cad63a;
sos_loop[0].somModel.tcam_mask[5][182][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][183][0]=80'h0000000016398c9c5329;
sos_loop[0].somModel.tcam_mask[5][183][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][184][0]=80'h00000000c1d9c5b84501;
sos_loop[0].somModel.tcam_mask[5][184][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][185][0]=80'h00000000d1ad3332662b;
sos_loop[0].somModel.tcam_mask[5][185][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][186][0]=80'h00000000b91d094ca5fa;
sos_loop[0].somModel.tcam_mask[5][186][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][187][0]=80'h0000000066807169ce5b;
sos_loop[0].somModel.tcam_mask[5][187][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][188][0]=80'h000000006ef096e4f564;
sos_loop[0].somModel.tcam_mask[5][188][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][189][0]=80'h00000000328864e675f7;
sos_loop[0].somModel.tcam_mask[5][189][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][190][0]=80'h000000007dae2b0e1b45;
sos_loop[0].somModel.tcam_mask[5][190][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][191][0]=80'h00000000bcb94b47b6e1;
sos_loop[0].somModel.tcam_mask[5][191][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][192][0]=80'h00000000969630df4be5;
sos_loop[0].somModel.tcam_mask[5][192][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][193][0]=80'h000000008fa1021a531a;
sos_loop[0].somModel.tcam_mask[5][193][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][194][0]=80'h00000000872d61d5debf;
sos_loop[0].somModel.tcam_mask[5][194][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][195][0]=80'h00000000991610788933;
sos_loop[0].somModel.tcam_mask[5][195][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][196][0]=80'h000000000abf899e0a35;
sos_loop[0].somModel.tcam_mask[5][196][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][197][0]=80'h000000009a50b37b4c4e;
sos_loop[0].somModel.tcam_mask[5][197][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][198][0]=80'h00000000a57859f9c477;
sos_loop[0].somModel.tcam_mask[5][198][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][199][0]=80'h000000000079cd60c49c;
sos_loop[0].somModel.tcam_mask[5][199][0]=80'hffffffffff8000000000;
sos_loop[0].somModel.tcam_data[5][200][0]=80'h00000000116a5a1abd7d;
sos_loop[0].somModel.tcam_mask[5][200][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][201][0]=80'h00000000c21fd0b46818;
sos_loop[0].somModel.tcam_mask[5][201][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][202][0]=80'h00000000cb7c1d8cfffa;
sos_loop[0].somModel.tcam_mask[5][202][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][203][0]=80'h000000005da2668e789f;
sos_loop[0].somModel.tcam_mask[5][203][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][204][0]=80'h00000000a975554d1660;
sos_loop[0].somModel.tcam_mask[5][204][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][205][0]=80'h00000000f527f8412a24;
sos_loop[0].somModel.tcam_mask[5][205][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][206][0]=80'h000000006e7cabe12a47;
sos_loop[0].somModel.tcam_mask[5][206][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][207][0]=80'h00000000ecce1c4cd86e;
sos_loop[0].somModel.tcam_mask[5][207][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][208][0]=80'h0000000072d3d3fcd72b;
sos_loop[0].somModel.tcam_mask[5][208][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][209][0]=80'h00000000839e1fb55d44;
sos_loop[0].somModel.tcam_mask[5][209][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][210][0]=80'h00000000478398e0b9ee;
sos_loop[0].somModel.tcam_mask[5][210][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][211][0]=80'h000000008530d50e759f;
sos_loop[0].somModel.tcam_mask[5][211][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][212][0]=80'h0000000011f968361ebd;
sos_loop[0].somModel.tcam_mask[5][212][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][213][0]=80'h000000008ce994cc083f;
sos_loop[0].somModel.tcam_mask[5][213][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][214][0]=80'h000000002c23f84988ee;
sos_loop[0].somModel.tcam_mask[5][214][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][215][0]=80'h000000009760938f25c2;
sos_loop[0].somModel.tcam_mask[5][215][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][216][0]=80'h00000000274efbfa8211;
sos_loop[0].somModel.tcam_mask[5][216][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][217][0]=80'h00000000694132b93ba3;
sos_loop[0].somModel.tcam_mask[5][217][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][218][0]=80'h000000000682f3056401;
sos_loop[0].somModel.tcam_mask[5][218][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][219][0]=80'h00000000d1c36a785d4f;
sos_loop[0].somModel.tcam_mask[5][219][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][220][0]=80'h000000004ae9b6d2ef4f;
sos_loop[0].somModel.tcam_mask[5][220][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][221][0]=80'h00000000c9c32ab41eeb;
sos_loop[0].somModel.tcam_mask[5][221][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][222][0]=80'h00000000cbc076ebe28e;
sos_loop[0].somModel.tcam_mask[5][222][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][223][0]=80'h00000000fbda31fd76c0;
sos_loop[0].somModel.tcam_mask[5][223][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][224][0]=80'h000000009a099a151b35;
sos_loop[0].somModel.tcam_mask[5][224][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][225][0]=80'h0000000054a1681b3ffb;
sos_loop[0].somModel.tcam_mask[5][225][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][226][0]=80'h00000000f0cf8f9ee272;
sos_loop[0].somModel.tcam_mask[5][226][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][227][0]=80'h000000003f535b44d28a;
sos_loop[0].somModel.tcam_mask[5][227][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][228][0]=80'h000000007ae44fa333c8;
sos_loop[0].somModel.tcam_mask[5][228][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][229][0]=80'h00000000b665ce7f735a;
sos_loop[0].somModel.tcam_mask[5][229][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][230][0]=80'h00000000626c7ae8774d;
sos_loop[0].somModel.tcam_mask[5][230][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][231][0]=80'h00000000f3cddb51d392;
sos_loop[0].somModel.tcam_mask[5][231][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][232][0]=80'h00000000944a75a8319c;
sos_loop[0].somModel.tcam_mask[5][232][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][233][0]=80'h00000000eaacb9890fae;
sos_loop[0].somModel.tcam_mask[5][233][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][234][0]=80'h00000000046f6540ec7f;
sos_loop[0].somModel.tcam_mask[5][234][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][235][0]=80'h00000000c6088fc1bd3d;
sos_loop[0].somModel.tcam_mask[5][235][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][236][0]=80'h000000005e0b61c56031;
sos_loop[0].somModel.tcam_mask[5][236][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][237][0]=80'h00000000027b4c51c3bb;
sos_loop[0].somModel.tcam_mask[5][237][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[5][238][0]=80'h00000000be4d82d7e60e;
sos_loop[0].somModel.tcam_mask[5][238][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][239][0]=80'h000000007eef6a0932c5;
sos_loop[0].somModel.tcam_mask[5][239][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][240][0]=80'h00000000564f40cb3bc6;
sos_loop[0].somModel.tcam_mask[5][240][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][241][0]=80'h0000000049ba0e14ede1;
sos_loop[0].somModel.tcam_mask[5][241][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][242][0]=80'h000000000ffa1385e8e1;
sos_loop[0].somModel.tcam_mask[5][242][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][243][0]=80'h00000000c2a6a6c5875c;
sos_loop[0].somModel.tcam_mask[5][243][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][244][0]=80'h0000000046ed88992ff9;
sos_loop[0].somModel.tcam_mask[5][244][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][245][0]=80'h000000007bd52c488741;
sos_loop[0].somModel.tcam_mask[5][245][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][246][0]=80'h00000000dd037b320186;
sos_loop[0].somModel.tcam_mask[5][246][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][247][0]=80'h00000000bc45bae8ac0a;
sos_loop[0].somModel.tcam_mask[5][247][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][248][0]=80'h000000005b06c7e96f30;
sos_loop[0].somModel.tcam_mask[5][248][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][249][0]=80'h00000000d4ddc557a673;
sos_loop[0].somModel.tcam_mask[5][249][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][250][0]=80'h0000000053ec21af6aa7;
sos_loop[0].somModel.tcam_mask[5][250][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][251][0]=80'h0000000017ac57f88e87;
sos_loop[0].somModel.tcam_mask[5][251][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][252][0]=80'h00000000a4100e4032cc;
sos_loop[0].somModel.tcam_mask[5][252][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][253][0]=80'h00000000140fa51dda60;
sos_loop[0].somModel.tcam_mask[5][253][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][254][0]=80'h00000000ba76b63b04af;
sos_loop[0].somModel.tcam_mask[5][254][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][255][0]=80'h000000007bf30212d42d;
sos_loop[0].somModel.tcam_mask[5][255][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][256][0]=80'h00000000389a856d0929;
sos_loop[0].somModel.tcam_mask[5][256][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][257][0]=80'h00000000971def77bfa0;
sos_loop[0].somModel.tcam_mask[5][257][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][258][0]=80'h000000007fea6ca2dda9;
sos_loop[0].somModel.tcam_mask[5][258][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][259][0]=80'h000000006cc87b7163e1;
sos_loop[0].somModel.tcam_mask[5][259][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][260][0]=80'h00000000652f37432033;
sos_loop[0].somModel.tcam_mask[5][260][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][261][0]=80'h0000000094ca0afeaf40;
sos_loop[0].somModel.tcam_mask[5][261][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][262][0]=80'h00000000aa6075a82cfd;
sos_loop[0].somModel.tcam_mask[5][262][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][263][0]=80'h00000000e393132fbd4d;
sos_loop[0].somModel.tcam_mask[5][263][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][264][0]=80'h000000008617fb8769a3;
sos_loop[0].somModel.tcam_mask[5][264][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][265][0]=80'h00000000d45704f554fa;
sos_loop[0].somModel.tcam_mask[5][265][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][266][0]=80'h00000000083aeac67707;
sos_loop[0].somModel.tcam_mask[5][266][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][267][0]=80'h00000000ad11dd592c9a;
sos_loop[0].somModel.tcam_mask[5][267][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][268][0]=80'h00000000199fcd09ed28;
sos_loop[0].somModel.tcam_mask[5][268][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][269][0]=80'h00000000306fc67d4fd2;
sos_loop[0].somModel.tcam_mask[5][269][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][270][0]=80'h00000000ded308236673;
sos_loop[0].somModel.tcam_mask[5][270][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][271][0]=80'h000000006bb4f3981543;
sos_loop[0].somModel.tcam_mask[5][271][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][272][0]=80'h0000000028d774fa8bab;
sos_loop[0].somModel.tcam_mask[5][272][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][273][0]=80'h000000005f39e126fa40;
sos_loop[0].somModel.tcam_mask[5][273][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][274][0]=80'h000000004ec1930dd830;
sos_loop[0].somModel.tcam_mask[5][274][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][275][0]=80'h000000002eabafa47444;
sos_loop[0].somModel.tcam_mask[5][275][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][276][0]=80'h00000000f2c4354979b5;
sos_loop[0].somModel.tcam_mask[5][276][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][277][0]=80'h000000004375ff2839ff;
sos_loop[0].somModel.tcam_mask[5][277][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][278][0]=80'h00000000831847d750e3;
sos_loop[0].somModel.tcam_mask[5][278][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][279][0]=80'h000000006d4ff70a7fc3;
sos_loop[0].somModel.tcam_mask[5][279][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][280][0]=80'h0000000067633ad96690;
sos_loop[0].somModel.tcam_mask[5][280][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][281][0]=80'h0000000058b1bb7ab35b;
sos_loop[0].somModel.tcam_mask[5][281][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][282][0]=80'h00000000378d65b1297a;
sos_loop[0].somModel.tcam_mask[5][282][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][283][0]=80'h000000008ab24a720a34;
sos_loop[0].somModel.tcam_mask[5][283][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][284][0]=80'h000000009b617faf808a;
sos_loop[0].somModel.tcam_mask[5][284][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][285][0]=80'h000000002b5be33345f9;
sos_loop[0].somModel.tcam_mask[5][285][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][286][0]=80'h0000000080b069925240;
sos_loop[0].somModel.tcam_mask[5][286][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][287][0]=80'h0000000064819ae5ce38;
sos_loop[0].somModel.tcam_mask[5][287][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][288][0]=80'h00000000c8a2886319ad;
sos_loop[0].somModel.tcam_mask[5][288][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][289][0]=80'h00000000bba80680cd74;
sos_loop[0].somModel.tcam_mask[5][289][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][290][0]=80'h00000000c624c1780420;
sos_loop[0].somModel.tcam_mask[5][290][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][291][0]=80'h000000000df4dc19f8a0;
sos_loop[0].somModel.tcam_mask[5][291][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][292][0]=80'h00000000bf4fc4c5109d;
sos_loop[0].somModel.tcam_mask[5][292][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][293][0]=80'h00000000230e53a6e40d;
sos_loop[0].somModel.tcam_mask[5][293][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][294][0]=80'h000000006a8845704812;
sos_loop[0].somModel.tcam_mask[5][294][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][295][0]=80'h00000000d02d7e61c3ff;
sos_loop[0].somModel.tcam_mask[5][295][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][296][0]=80'h0000000042d9ad4b7cb5;
sos_loop[0].somModel.tcam_mask[5][296][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][297][0]=80'h000000006620c43e40cd;
sos_loop[0].somModel.tcam_mask[5][297][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][298][0]=80'h00000000572b2a5075a9;
sos_loop[0].somModel.tcam_mask[5][298][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][299][0]=80'h000000000bc0a3cd8632;
sos_loop[0].somModel.tcam_mask[5][299][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][300][0]=80'h00000000318840f45c23;
sos_loop[0].somModel.tcam_mask[5][300][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][301][0]=80'h000000007ec0b9f2df84;
sos_loop[0].somModel.tcam_mask[5][301][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][302][0]=80'h000000000708eaeea371;
sos_loop[0].somModel.tcam_mask[5][302][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][303][0]=80'h0000000029e3e9901c1f;
sos_loop[0].somModel.tcam_mask[5][303][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][304][0]=80'h00000000f4f0fb40376f;
sos_loop[0].somModel.tcam_mask[5][304][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][305][0]=80'h000000007de8c27c7bf8;
sos_loop[0].somModel.tcam_mask[5][305][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][306][0]=80'h00000000722214538bb3;
sos_loop[0].somModel.tcam_mask[5][306][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][307][0]=80'h00000000b35284a2e8f3;
sos_loop[0].somModel.tcam_mask[5][307][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][308][0]=80'h00000000c1e963dc4088;
sos_loop[0].somModel.tcam_mask[5][308][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][309][0]=80'h0000000050d5503770e6;
sos_loop[0].somModel.tcam_mask[5][309][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][310][0]=80'h00000000b63951662a30;
sos_loop[0].somModel.tcam_mask[5][310][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][311][0]=80'h000000007eddea567619;
sos_loop[0].somModel.tcam_mask[5][311][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][312][0]=80'h000000004eab0a109e8f;
sos_loop[0].somModel.tcam_mask[5][312][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][313][0]=80'h00000000e549f26a551a;
sos_loop[0].somModel.tcam_mask[5][313][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][314][0]=80'h00000000161e12d7d5f4;
sos_loop[0].somModel.tcam_mask[5][314][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][315][0]=80'h000000002fb8691cf03d;
sos_loop[0].somModel.tcam_mask[5][315][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][316][0]=80'h000000006d0dd414bd88;
sos_loop[0].somModel.tcam_mask[5][316][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][317][0]=80'h00000000d47f0cfd8269;
sos_loop[0].somModel.tcam_mask[5][317][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][318][0]=80'h00000000e7fe58f76aac;
sos_loop[0].somModel.tcam_mask[5][318][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][319][0]=80'h00000000cddb5437e4b9;
sos_loop[0].somModel.tcam_mask[5][319][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][320][0]=80'h0000000058ac2d7d65c1;
sos_loop[0].somModel.tcam_mask[5][320][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][321][0]=80'h00000000e81d8eb85034;
sos_loop[0].somModel.tcam_mask[5][321][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][322][0]=80'h00000000a6fb99d69d1b;
sos_loop[0].somModel.tcam_mask[5][322][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][323][0]=80'h0000000085db0f2ad52e;
sos_loop[0].somModel.tcam_mask[5][323][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][324][0]=80'h00000000ba447f49c0b1;
sos_loop[0].somModel.tcam_mask[5][324][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][325][0]=80'h0000000099d3496acd35;
sos_loop[0].somModel.tcam_mask[5][325][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][326][0]=80'h0000000040e7e1b07303;
sos_loop[0].somModel.tcam_mask[5][326][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][327][0]=80'h0000000055f948ebe91d;
sos_loop[0].somModel.tcam_mask[5][327][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][328][0]=80'h00000000392c0459ce02;
sos_loop[0].somModel.tcam_mask[5][328][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][329][0]=80'h000000007e3d419f5d34;
sos_loop[0].somModel.tcam_mask[5][329][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][330][0]=80'h00000000e74efb58eaa7;
sos_loop[0].somModel.tcam_mask[5][330][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][331][0]=80'h00000000f83f581e4482;
sos_loop[0].somModel.tcam_mask[5][331][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][332][0]=80'h000000009cce1dfeef14;
sos_loop[0].somModel.tcam_mask[5][332][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][333][0]=80'h000000004b70936e9f64;
sos_loop[0].somModel.tcam_mask[5][333][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][334][0]=80'h000000008f60bf446783;
sos_loop[0].somModel.tcam_mask[5][334][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][335][0]=80'h0000000093a9046448e2;
sos_loop[0].somModel.tcam_mask[5][335][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][336][0]=80'h000000006e3ce4ac6730;
sos_loop[0].somModel.tcam_mask[5][336][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][337][0]=80'h0000000084de22fbc40a;
sos_loop[0].somModel.tcam_mask[5][337][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][338][0]=80'h000000002d98732c0914;
sos_loop[0].somModel.tcam_mask[5][338][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][339][0]=80'h00000000588e0584287c;
sos_loop[0].somModel.tcam_mask[5][339][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][340][0]=80'h000000008f50e0497e89;
sos_loop[0].somModel.tcam_mask[5][340][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][341][0]=80'h00000000b0e119fb2555;
sos_loop[0].somModel.tcam_mask[5][341][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][342][0]=80'h000000004cd3c2cde21a;
sos_loop[0].somModel.tcam_mask[5][342][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][343][0]=80'h00000000da342cb3beee;
sos_loop[0].somModel.tcam_mask[5][343][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][344][0]=80'h000000009f7fc5e6a042;
sos_loop[0].somModel.tcam_mask[5][344][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][345][0]=80'h00000000cc5300c82669;
sos_loop[0].somModel.tcam_mask[5][345][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][346][0]=80'h000000006a1ec386bf00;
sos_loop[0].somModel.tcam_mask[5][346][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][347][0]=80'h000000002317e8d90545;
sos_loop[0].somModel.tcam_mask[5][347][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][348][0]=80'h000000008d4fe98625cf;
sos_loop[0].somModel.tcam_mask[5][348][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][349][0]=80'h00000000060665e2c19e;
sos_loop[0].somModel.tcam_mask[5][349][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][350][0]=80'h00000000596674fbbfb1;
sos_loop[0].somModel.tcam_mask[5][350][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][351][0]=80'h000000005c7688d8aad5;
sos_loop[0].somModel.tcam_mask[5][351][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][352][0]=80'h0000000099c3cb202d30;
sos_loop[0].somModel.tcam_mask[5][352][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][353][0]=80'h00000000a86ac83a7681;
sos_loop[0].somModel.tcam_mask[5][353][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][354][0]=80'h00000000f9f330aaf7e5;
sos_loop[0].somModel.tcam_mask[5][354][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][355][0]=80'h000000003c3dcdb988e5;
sos_loop[0].somModel.tcam_mask[5][355][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][356][0]=80'h0000000082440e73e0a4;
sos_loop[0].somModel.tcam_mask[5][356][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][357][0]=80'h00000000deb63d376bdd;
sos_loop[0].somModel.tcam_mask[5][357][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][358][0]=80'h000000003f13c6d986da;
sos_loop[0].somModel.tcam_mask[5][358][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][359][0]=80'h00000000959a11161a8a;
sos_loop[0].somModel.tcam_mask[5][359][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][360][0]=80'h0000000004fc4b9709a2;
sos_loop[0].somModel.tcam_mask[5][360][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][361][0]=80'h000000000603260a4fa8;
sos_loop[0].somModel.tcam_mask[5][361][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][362][0]=80'h00000000317642426d30;
sos_loop[0].somModel.tcam_mask[5][362][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][363][0]=80'h0000000093eea5159da0;
sos_loop[0].somModel.tcam_mask[5][363][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][364][0]=80'h00000000a6a6c5effbb8;
sos_loop[0].somModel.tcam_mask[5][364][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][365][0]=80'h000000009a556fc0f1e1;
sos_loop[0].somModel.tcam_mask[5][365][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][366][0]=80'h00000000ca8bfde422b1;
sos_loop[0].somModel.tcam_mask[5][366][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][367][0]=80'h000000006b3d4da4a0e4;
sos_loop[0].somModel.tcam_mask[5][367][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][368][0]=80'h00000000b8725432eee0;
sos_loop[0].somModel.tcam_mask[5][368][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][369][0]=80'h000000002a5f4d97572c;
sos_loop[0].somModel.tcam_mask[5][369][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][370][0]=80'h0000000003f4b2f37c91;
sos_loop[0].somModel.tcam_mask[5][370][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[5][371][0]=80'h000000006d012a56f306;
sos_loop[0].somModel.tcam_mask[5][371][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][372][0]=80'h00000000f39c18ff7423;
sos_loop[0].somModel.tcam_mask[5][372][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][373][0]=80'h0000000064fe54c3d020;
sos_loop[0].somModel.tcam_mask[5][373][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][374][0]=80'h000000005941386df853;
sos_loop[0].somModel.tcam_mask[5][374][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][375][0]=80'h00000000fd5081a7023d;
sos_loop[0].somModel.tcam_mask[5][375][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][376][0]=80'h0000000059d252677e44;
sos_loop[0].somModel.tcam_mask[5][376][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][377][0]=80'h00000000b1ef710456c8;
sos_loop[0].somModel.tcam_mask[5][377][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][378][0]=80'h000000008a3b29afa55f;
sos_loop[0].somModel.tcam_mask[5][378][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][379][0]=80'h00000000a8f4af7c920a;
sos_loop[0].somModel.tcam_mask[5][379][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][380][0]=80'h000000009b5b556528f0;
sos_loop[0].somModel.tcam_mask[5][380][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][381][0]=80'h000000008d75c4ce6384;
sos_loop[0].somModel.tcam_mask[5][381][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][382][0]=80'h00000000644e172a4d39;
sos_loop[0].somModel.tcam_mask[5][382][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][383][0]=80'h000000004e2c31c4e9bf;
sos_loop[0].somModel.tcam_mask[5][383][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][384][0]=80'h00000000fb16e104670e;
sos_loop[0].somModel.tcam_mask[5][384][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][385][0]=80'h00000000edda66338267;
sos_loop[0].somModel.tcam_mask[5][385][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][386][0]=80'h00000000028c12a16f1b;
sos_loop[0].somModel.tcam_mask[5][386][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[5][387][0]=80'h00000000ff84824ad314;
sos_loop[0].somModel.tcam_mask[5][387][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][388][0]=80'h000000000be7756aeeab;
sos_loop[0].somModel.tcam_mask[5][388][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][389][0]=80'h000000007e61e055303f;
sos_loop[0].somModel.tcam_mask[5][389][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][390][0]=80'h00000000aac7193a22af;
sos_loop[0].somModel.tcam_mask[5][390][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][391][0]=80'h00000000565f0106873e;
sos_loop[0].somModel.tcam_mask[5][391][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][392][0]=80'h0000000075032e61802d;
sos_loop[0].somModel.tcam_mask[5][392][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][393][0]=80'h00000000f2f7c9dbbf6e;
sos_loop[0].somModel.tcam_mask[5][393][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][394][0]=80'h00000000c616b82074dc;
sos_loop[0].somModel.tcam_mask[5][394][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][395][0]=80'h000000009b90c73a26b9;
sos_loop[0].somModel.tcam_mask[5][395][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][396][0]=80'h00000000f1aad48501e0;
sos_loop[0].somModel.tcam_mask[5][396][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][397][0]=80'h00000000b50e5a5b2331;
sos_loop[0].somModel.tcam_mask[5][397][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][398][0]=80'h000000000536e70ff511;
sos_loop[0].somModel.tcam_mask[5][398][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][399][0]=80'h00000000500f137223d6;
sos_loop[0].somModel.tcam_mask[5][399][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][400][0]=80'h000000002791051b62a6;
sos_loop[0].somModel.tcam_mask[5][400][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][401][0]=80'h00000000c4eb2c045df0;
sos_loop[0].somModel.tcam_mask[5][401][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][402][0]=80'h00000000a4ad1b4e4c65;
sos_loop[0].somModel.tcam_mask[5][402][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][403][0]=80'h000000005dcd203c62ab;
sos_loop[0].somModel.tcam_mask[5][403][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][404][0]=80'h00000000bd2053fe1aa1;
sos_loop[0].somModel.tcam_mask[5][404][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][405][0]=80'h00000000dd873733eebd;
sos_loop[0].somModel.tcam_mask[5][405][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][406][0]=80'h00000000d5cc8944cc44;
sos_loop[0].somModel.tcam_mask[5][406][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][407][0]=80'h00000000df75e34c1d60;
sos_loop[0].somModel.tcam_mask[5][407][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][408][0]=80'h0000000069516c90e02b;
sos_loop[0].somModel.tcam_mask[5][408][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][409][0]=80'h00000000ba7434218648;
sos_loop[0].somModel.tcam_mask[5][409][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][410][0]=80'h0000000075995e082cc9;
sos_loop[0].somModel.tcam_mask[5][410][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][411][0]=80'h000000008f8a0618c492;
sos_loop[0].somModel.tcam_mask[5][411][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][412][0]=80'h0000000085652adefb50;
sos_loop[0].somModel.tcam_mask[5][412][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][413][0]=80'h0000000084e3bbb346a9;
sos_loop[0].somModel.tcam_mask[5][413][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][414][0]=80'h00000000ce288545ff5c;
sos_loop[0].somModel.tcam_mask[5][414][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][415][0]=80'h00000000f34840529bc7;
sos_loop[0].somModel.tcam_mask[5][415][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][416][0]=80'h0000000093b680734ca8;
sos_loop[0].somModel.tcam_mask[5][416][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][417][0]=80'h000000006d3e5930bf31;
sos_loop[0].somModel.tcam_mask[5][417][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][418][0]=80'h000000004c6bb4e13dd2;
sos_loop[0].somModel.tcam_mask[5][418][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][419][0]=80'h00000000c17e7cae146d;
sos_loop[0].somModel.tcam_mask[5][419][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][420][0]=80'h000000003a01e234f448;
sos_loop[0].somModel.tcam_mask[5][420][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][421][0]=80'h000000001f6089a70d31;
sos_loop[0].somModel.tcam_mask[5][421][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][422][0]=80'h00000000e9910acedf01;
sos_loop[0].somModel.tcam_mask[5][422][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][423][0]=80'h0000000092c1be63a45c;
sos_loop[0].somModel.tcam_mask[5][423][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][424][0]=80'h0000000077250b5545e8;
sos_loop[0].somModel.tcam_mask[5][424][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][425][0]=80'h0000000041875a4af1b4;
sos_loop[0].somModel.tcam_mask[5][425][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][426][0]=80'h000000001f7188b8f195;
sos_loop[0].somModel.tcam_mask[5][426][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][427][0]=80'h00000000e7043697f5e9;
sos_loop[0].somModel.tcam_mask[5][427][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][428][0]=80'h00000000ccb0a5325cbe;
sos_loop[0].somModel.tcam_mask[5][428][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][429][0]=80'h00000000f77c99d0ae10;
sos_loop[0].somModel.tcam_mask[5][429][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][430][0]=80'h0000000051c66267cec7;
sos_loop[0].somModel.tcam_mask[5][430][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][431][0]=80'h00000000a3eb7b517f7d;
sos_loop[0].somModel.tcam_mask[5][431][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][432][0]=80'h000000005e4b84a9a324;
sos_loop[0].somModel.tcam_mask[5][432][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][433][0]=80'h00000000263366d9a934;
sos_loop[0].somModel.tcam_mask[5][433][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][434][0]=80'h0000000035cd167e2bad;
sos_loop[0].somModel.tcam_mask[5][434][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][435][0]=80'h000000000b2c3bbf8fba;
sos_loop[0].somModel.tcam_mask[5][435][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][436][0]=80'h000000008f19a66976c7;
sos_loop[0].somModel.tcam_mask[5][436][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][437][0]=80'h00000000e0b42c35622b;
sos_loop[0].somModel.tcam_mask[5][437][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][438][0]=80'h00000000dca9a6f1782c;
sos_loop[0].somModel.tcam_mask[5][438][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][439][0]=80'h000000009a1541c274a2;
sos_loop[0].somModel.tcam_mask[5][439][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][440][0]=80'h0000000044768a38b95d;
sos_loop[0].somModel.tcam_mask[5][440][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][441][0]=80'h0000000038f48a68b142;
sos_loop[0].somModel.tcam_mask[5][441][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][442][0]=80'h000000009759c188b4fd;
sos_loop[0].somModel.tcam_mask[5][442][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][443][0]=80'h00000000a08c0f3399b6;
sos_loop[0].somModel.tcam_mask[5][443][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][444][0]=80'h00000000820dea118ef9;
sos_loop[0].somModel.tcam_mask[5][444][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][445][0]=80'h00000000786f4fec3569;
sos_loop[0].somModel.tcam_mask[5][445][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][446][0]=80'h0000000035502a9bf339;
sos_loop[0].somModel.tcam_mask[5][446][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][447][0]=80'h00000000ede032f81911;
sos_loop[0].somModel.tcam_mask[5][447][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][448][0]=80'h00000000005d2da41d57;
sos_loop[0].somModel.tcam_mask[5][448][0]=80'hffffffffff8000000000;
sos_loop[0].somModel.tcam_data[5][449][0]=80'h000000001d551e45233a;
sos_loop[0].somModel.tcam_mask[5][449][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][450][0]=80'h000000001232e7e21619;
sos_loop[0].somModel.tcam_mask[5][450][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][451][0]=80'h000000009656bf8e0b9d;
sos_loop[0].somModel.tcam_mask[5][451][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][452][0]=80'h00000000282df63c9a42;
sos_loop[0].somModel.tcam_mask[5][452][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][453][0]=80'h00000000fb8cfa3efc1a;
sos_loop[0].somModel.tcam_mask[5][453][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][454][0]=80'h00000000e202a5e04142;
sos_loop[0].somModel.tcam_mask[5][454][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][455][0]=80'h00000000ce14bd93ed55;
sos_loop[0].somModel.tcam_mask[5][455][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][456][0]=80'h000000000b29b6b75332;
sos_loop[0].somModel.tcam_mask[5][456][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][457][0]=80'h00000000a560cfe7acfc;
sos_loop[0].somModel.tcam_mask[5][457][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][458][0]=80'h0000000099c7f0448e01;
sos_loop[0].somModel.tcam_mask[5][458][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][459][0]=80'h000000001dc007e9c85a;
sos_loop[0].somModel.tcam_mask[5][459][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][460][0]=80'h00000000d5bbfcebded1;
sos_loop[0].somModel.tcam_mask[5][460][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][461][0]=80'h000000007a59ce859cc7;
sos_loop[0].somModel.tcam_mask[5][461][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][462][0]=80'h000000004ea8c5b70bda;
sos_loop[0].somModel.tcam_mask[5][462][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][463][0]=80'h0000000052f1807fc08a;
sos_loop[0].somModel.tcam_mask[5][463][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][464][0]=80'h00000000206171d9529a;
sos_loop[0].somModel.tcam_mask[5][464][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][465][0]=80'h00000000498a7ea9d6a4;
sos_loop[0].somModel.tcam_mask[5][465][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][466][0]=80'h0000000068b1d8990008;
sos_loop[0].somModel.tcam_mask[5][466][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][467][0]=80'h00000000dfdd7f5c6649;
sos_loop[0].somModel.tcam_mask[5][467][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][468][0]=80'h00000000423c83f43d47;
sos_loop[0].somModel.tcam_mask[5][468][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][469][0]=80'h0000000071daa74440c3;
sos_loop[0].somModel.tcam_mask[5][469][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][470][0]=80'h000000006b7caeb2cb69;
sos_loop[0].somModel.tcam_mask[5][470][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][471][0]=80'h000000009301716b199f;
sos_loop[0].somModel.tcam_mask[5][471][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][472][0]=80'h00000000f30c2c261355;
sos_loop[0].somModel.tcam_mask[5][472][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][473][0]=80'h00000000e1037b5789b6;
sos_loop[0].somModel.tcam_mask[5][473][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][474][0]=80'h000000004ac85c163c30;
sos_loop[0].somModel.tcam_mask[5][474][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][475][0]=80'h00000000bd2e17a3bd71;
sos_loop[0].somModel.tcam_mask[5][475][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][476][0]=80'h000000008cfbaac12a25;
sos_loop[0].somModel.tcam_mask[5][476][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][477][0]=80'h00000000e07f86b355a4;
sos_loop[0].somModel.tcam_mask[5][477][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][478][0]=80'h00000000e24b3b5f435d;
sos_loop[0].somModel.tcam_mask[5][478][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][479][0]=80'h00000000c6100a3221e3;
sos_loop[0].somModel.tcam_mask[5][479][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][480][0]=80'h00000000d601e9e5d6ac;
sos_loop[0].somModel.tcam_mask[5][480][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][481][0]=80'h00000000a2ee82f9007b;
sos_loop[0].somModel.tcam_mask[5][481][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][482][0]=80'h00000000b4baf8944204;
sos_loop[0].somModel.tcam_mask[5][482][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][483][0]=80'h0000000078c5ee1f506d;
sos_loop[0].somModel.tcam_mask[5][483][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][484][0]=80'h0000000094176a64d950;
sos_loop[0].somModel.tcam_mask[5][484][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][485][0]=80'h00000000bdc7edf2bed3;
sos_loop[0].somModel.tcam_mask[5][485][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][486][0]=80'h00000000f6141087125a;
sos_loop[0].somModel.tcam_mask[5][486][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][487][0]=80'h000000004d8a6c4bb175;
sos_loop[0].somModel.tcam_mask[5][487][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][488][0]=80'h00000000d702b7ff755e;
sos_loop[0].somModel.tcam_mask[5][488][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][489][0]=80'h0000000017ad459c4491;
sos_loop[0].somModel.tcam_mask[5][489][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][490][0]=80'h00000000becd69de0af5;
sos_loop[0].somModel.tcam_mask[5][490][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][491][0]=80'h000000006db83a09cb40;
sos_loop[0].somModel.tcam_mask[5][491][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][492][0]=80'h00000000c15a3192c54e;
sos_loop[0].somModel.tcam_mask[5][492][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][493][0]=80'h00000000372729de79a7;
sos_loop[0].somModel.tcam_mask[5][493][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][494][0]=80'h00000000b7d5a573112e;
sos_loop[0].somModel.tcam_mask[5][494][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][495][0]=80'h00000000e7598a8d64ef;
sos_loop[0].somModel.tcam_mask[5][495][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][496][0]=80'h000000004d77a8f186e8;
sos_loop[0].somModel.tcam_mask[5][496][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][497][0]=80'h00000000b3a7e8c62438;
sos_loop[0].somModel.tcam_mask[5][497][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][498][0]=80'h000000005e628e40bad8;
sos_loop[0].somModel.tcam_mask[5][498][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][499][0]=80'h000000002c6ae9566a81;
sos_loop[0].somModel.tcam_mask[5][499][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][500][0]=80'h000000007c8088a4d780;
sos_loop[0].somModel.tcam_mask[5][500][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][501][0]=80'h00000000449da718991b;
sos_loop[0].somModel.tcam_mask[5][501][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][502][0]=80'h00000000eb14915c851e;
sos_loop[0].somModel.tcam_mask[5][502][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][503][0]=80'h000000003527b3d245b5;
sos_loop[0].somModel.tcam_mask[5][503][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][504][0]=80'h0000000085d7cc131a8a;
sos_loop[0].somModel.tcam_mask[5][504][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][505][0]=80'h00000000b448dcc734b3;
sos_loop[0].somModel.tcam_mask[5][505][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][506][0]=80'h000000000463282aaf56;
sos_loop[0].somModel.tcam_mask[5][506][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][507][0]=80'h00000000e6f6fe35b667;
sos_loop[0].somModel.tcam_mask[5][507][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][508][0]=80'h0000000080c258b15826;
sos_loop[0].somModel.tcam_mask[5][508][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][509][0]=80'h00000000faac4f7283f1;
sos_loop[0].somModel.tcam_mask[5][509][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][510][0]=80'h00000000a03cce697a88;
sos_loop[0].somModel.tcam_mask[5][510][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][511][0]=80'h00000000df03c7e186d0;
sos_loop[0].somModel.tcam_mask[5][511][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][512][0]=80'h00000000c301b2ddb491;
sos_loop[0].somModel.tcam_mask[5][512][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][513][0]=80'h0000000005a553a6d946;
sos_loop[0].somModel.tcam_mask[5][513][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][514][0]=80'h00000000ec81a0ecf565;
sos_loop[0].somModel.tcam_mask[5][514][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][515][0]=80'h0000000025b7ba6c7a22;
sos_loop[0].somModel.tcam_mask[5][515][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][516][0]=80'h00000000ff62f77af68e;
sos_loop[0].somModel.tcam_mask[5][516][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][517][0]=80'h0000000090696c0e7c49;
sos_loop[0].somModel.tcam_mask[5][517][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][518][0]=80'h00000000db542752b51b;
sos_loop[0].somModel.tcam_mask[5][518][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][519][0]=80'h000000005c669d7e5719;
sos_loop[0].somModel.tcam_mask[5][519][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][520][0]=80'h0000000007869b90d6d6;
sos_loop[0].somModel.tcam_mask[5][520][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][521][0]=80'h000000006ab3f4028bc4;
sos_loop[0].somModel.tcam_mask[5][521][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][522][0]=80'h00000000faf254c81784;
sos_loop[0].somModel.tcam_mask[5][522][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][523][0]=80'h00000000e91e80ddf2b6;
sos_loop[0].somModel.tcam_mask[5][523][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][524][0]=80'h0000000012ec8002dccf;
sos_loop[0].somModel.tcam_mask[5][524][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][525][0]=80'h000000001fb66119b301;
sos_loop[0].somModel.tcam_mask[5][525][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][526][0]=80'h0000000035cfa56dca6a;
sos_loop[0].somModel.tcam_mask[5][526][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][527][0]=80'h00000000257f17287640;
sos_loop[0].somModel.tcam_mask[5][527][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][528][0]=80'h00000000e24b719e5fd5;
sos_loop[0].somModel.tcam_mask[5][528][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][529][0]=80'h000000001b6de98d63bb;
sos_loop[0].somModel.tcam_mask[5][529][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][530][0]=80'h00000000c7396a1e1d0b;
sos_loop[0].somModel.tcam_mask[5][530][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][531][0]=80'h000000007fb43ae9cd4b;
sos_loop[0].somModel.tcam_mask[5][531][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][532][0]=80'h00000000a389a8825008;
sos_loop[0].somModel.tcam_mask[5][532][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][533][0]=80'h0000000062002cc089d3;
sos_loop[0].somModel.tcam_mask[5][533][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][534][0]=80'h00000000a2fc3e097fd8;
sos_loop[0].somModel.tcam_mask[5][534][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][535][0]=80'h0000000093938f2e7bb6;
sos_loop[0].somModel.tcam_mask[5][535][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][536][0]=80'h000000004c0878c8f3c9;
sos_loop[0].somModel.tcam_mask[5][536][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][537][0]=80'h000000006dad4681d74b;
sos_loop[0].somModel.tcam_mask[5][537][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][538][0]=80'h0000000090d849afd440;
sos_loop[0].somModel.tcam_mask[5][538][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][539][0]=80'h0000000099cea5c192b2;
sos_loop[0].somModel.tcam_mask[5][539][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][540][0]=80'h00000000439a63924ef9;
sos_loop[0].somModel.tcam_mask[5][540][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][541][0]=80'h0000000022efe4c3db4e;
sos_loop[0].somModel.tcam_mask[5][541][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][542][0]=80'h00000000935f8ae1eaca;
sos_loop[0].somModel.tcam_mask[5][542][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][543][0]=80'h00000000980ce89cb3ca;
sos_loop[0].somModel.tcam_mask[5][543][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][544][0]=80'h00000000b2b1d54e6143;
sos_loop[0].somModel.tcam_mask[5][544][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][545][0]=80'h00000000985262ca09c2;
sos_loop[0].somModel.tcam_mask[5][545][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][546][0]=80'h000000001b5370c23148;
sos_loop[0].somModel.tcam_mask[5][546][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][547][0]=80'h00000000fa6e44897737;
sos_loop[0].somModel.tcam_mask[5][547][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][548][0]=80'h00000000edc347b5f551;
sos_loop[0].somModel.tcam_mask[5][548][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][549][0]=80'h00000000bbafbcb86844;
sos_loop[0].somModel.tcam_mask[5][549][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][550][0]=80'h000000007fb9ba95cb59;
sos_loop[0].somModel.tcam_mask[5][550][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][551][0]=80'h00000000be931b35ee21;
sos_loop[0].somModel.tcam_mask[5][551][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][552][0]=80'h0000000039f56d709e34;
sos_loop[0].somModel.tcam_mask[5][552][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][553][0]=80'h000000004e9dfa08200a;
sos_loop[0].somModel.tcam_mask[5][553][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][554][0]=80'h00000000820c31b21a45;
sos_loop[0].somModel.tcam_mask[5][554][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][555][0]=80'h0000000005c7809f7005;
sos_loop[0].somModel.tcam_mask[5][555][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][556][0]=80'h000000003aca0c094cca;
sos_loop[0].somModel.tcam_mask[5][556][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][557][0]=80'h00000000745ae42f60b0;
sos_loop[0].somModel.tcam_mask[5][557][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][558][0]=80'h000000009ab1034e7c6e;
sos_loop[0].somModel.tcam_mask[5][558][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][559][0]=80'h000000008b03e00b02c2;
sos_loop[0].somModel.tcam_mask[5][559][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][560][0]=80'h00000000291393c268aa;
sos_loop[0].somModel.tcam_mask[5][560][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][561][0]=80'h000000004f5dda910b46;
sos_loop[0].somModel.tcam_mask[5][561][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][562][0]=80'h000000000d702572b740;
sos_loop[0].somModel.tcam_mask[5][562][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][563][0]=80'h0000000082eb751a50eb;
sos_loop[0].somModel.tcam_mask[5][563][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][564][0]=80'h0000000069f1bf212be5;
sos_loop[0].somModel.tcam_mask[5][564][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][565][0]=80'h00000000692f8eeae2e9;
sos_loop[0].somModel.tcam_mask[5][565][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][566][0]=80'h0000000019a683169415;
sos_loop[0].somModel.tcam_mask[5][566][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][567][0]=80'h0000000093bac3e6e685;
sos_loop[0].somModel.tcam_mask[5][567][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][568][0]=80'h000000004993bee769ac;
sos_loop[0].somModel.tcam_mask[5][568][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][569][0]=80'h00000000cd7fb4cb6753;
sos_loop[0].somModel.tcam_mask[5][569][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][570][0]=80'h000000000240e7a3c36d;
sos_loop[0].somModel.tcam_mask[5][570][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[5][571][0]=80'h00000000dee7cb29be85;
sos_loop[0].somModel.tcam_mask[5][571][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][572][0]=80'h00000000992597565e42;
sos_loop[0].somModel.tcam_mask[5][572][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][573][0]=80'h000000005cf48819c736;
sos_loop[0].somModel.tcam_mask[5][573][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][574][0]=80'h0000000047abe210da7f;
sos_loop[0].somModel.tcam_mask[5][574][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][575][0]=80'h00000000f93a1757baa0;
sos_loop[0].somModel.tcam_mask[5][575][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][576][0]=80'h000000007c1ceb4afc56;
sos_loop[0].somModel.tcam_mask[5][576][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][577][0]=80'h00000000af7d256d7cc4;
sos_loop[0].somModel.tcam_mask[5][577][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][578][0]=80'h0000000056f4eacb32c7;
sos_loop[0].somModel.tcam_mask[5][578][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][579][0]=80'h00000000b0d1add53e47;
sos_loop[0].somModel.tcam_mask[5][579][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][580][0]=80'h00000000d2755cc4bd17;
sos_loop[0].somModel.tcam_mask[5][580][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][581][0]=80'h00000000a6985589f9f2;
sos_loop[0].somModel.tcam_mask[5][581][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][582][0]=80'h00000000c617a79d7ece;
sos_loop[0].somModel.tcam_mask[5][582][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][583][0]=80'h00000000ce74602fffba;
sos_loop[0].somModel.tcam_mask[5][583][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][584][0]=80'h00000000f924b4b96d61;
sos_loop[0].somModel.tcam_mask[5][584][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][585][0]=80'h000000008c0b6b9901dc;
sos_loop[0].somModel.tcam_mask[5][585][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][586][0]=80'h00000000f68af87708bf;
sos_loop[0].somModel.tcam_mask[5][586][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][587][0]=80'h0000000074fa5f30fe3f;
sos_loop[0].somModel.tcam_mask[5][587][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][588][0]=80'h000000004db8a921b1d2;
sos_loop[0].somModel.tcam_mask[5][588][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][589][0]=80'h0000000018a72f979e24;
sos_loop[0].somModel.tcam_mask[5][589][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][590][0]=80'h00000000595e18260e26;
sos_loop[0].somModel.tcam_mask[5][590][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][591][0]=80'h00000000aad2d483e822;
sos_loop[0].somModel.tcam_mask[5][591][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][592][0]=80'h00000000343913fad305;
sos_loop[0].somModel.tcam_mask[5][592][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][593][0]=80'h00000000b3d2b6c10e97;
sos_loop[0].somModel.tcam_mask[5][593][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][594][0]=80'h000000005b359f4f70b0;
sos_loop[0].somModel.tcam_mask[5][594][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][595][0]=80'h00000000910fdf65238e;
sos_loop[0].somModel.tcam_mask[5][595][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][596][0]=80'h00000000858d2a03d342;
sos_loop[0].somModel.tcam_mask[5][596][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][597][0]=80'h0000000060c0b6079327;
sos_loop[0].somModel.tcam_mask[5][597][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][598][0]=80'h00000000ac7bf03559d7;
sos_loop[0].somModel.tcam_mask[5][598][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][599][0]=80'h000000009ad2390bbe32;
sos_loop[0].somModel.tcam_mask[5][599][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][600][0]=80'h00000000fa4f7ce06718;
sos_loop[0].somModel.tcam_mask[5][600][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][601][0]=80'h00000000d16fe65ec39f;
sos_loop[0].somModel.tcam_mask[5][601][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][602][0]=80'h000000002d99e55053a9;
sos_loop[0].somModel.tcam_mask[5][602][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][603][0]=80'h000000005159029f3697;
sos_loop[0].somModel.tcam_mask[5][603][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][604][0]=80'h00000000b4b0447b5549;
sos_loop[0].somModel.tcam_mask[5][604][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][605][0]=80'h00000000377b752a37b6;
sos_loop[0].somModel.tcam_mask[5][605][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][606][0]=80'h00000000220bb11437f4;
sos_loop[0].somModel.tcam_mask[5][606][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][607][0]=80'h00000000abd69fb1204e;
sos_loop[0].somModel.tcam_mask[5][607][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][608][0]=80'h00000000eb47988d0d8b;
sos_loop[0].somModel.tcam_mask[5][608][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][609][0]=80'h00000000ca9cc767edce;
sos_loop[0].somModel.tcam_mask[5][609][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][610][0]=80'h000000003b6f42cbe0a9;
sos_loop[0].somModel.tcam_mask[5][610][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][611][0]=80'h000000001dd3fa287076;
sos_loop[0].somModel.tcam_mask[5][611][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][612][0]=80'h000000009628912dbff2;
sos_loop[0].somModel.tcam_mask[5][612][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][613][0]=80'h0000000089a7951bea35;
sos_loop[0].somModel.tcam_mask[5][613][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][614][0]=80'h00000000c7b2ff90ab75;
sos_loop[0].somModel.tcam_mask[5][614][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][615][0]=80'h000000007ec37d3f35d1;
sos_loop[0].somModel.tcam_mask[5][615][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][616][0]=80'h00000000486d45350ba4;
sos_loop[0].somModel.tcam_mask[5][616][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][617][0]=80'h00000000f7c78a4aeffd;
sos_loop[0].somModel.tcam_mask[5][617][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][618][0]=80'h00000000ea7f3c4470a0;
sos_loop[0].somModel.tcam_mask[5][618][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][619][0]=80'h0000000095398bca46db;
sos_loop[0].somModel.tcam_mask[5][619][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][620][0]=80'h0000000002a21d269ef9;
sos_loop[0].somModel.tcam_mask[5][620][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[5][621][0]=80'h000000005ff142432afa;
sos_loop[0].somModel.tcam_mask[5][621][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][622][0]=80'h000000008d346fc65e2b;
sos_loop[0].somModel.tcam_mask[5][622][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][623][0]=80'h000000001a6584f50556;
sos_loop[0].somModel.tcam_mask[5][623][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][624][0]=80'h0000000008386da1029f;
sos_loop[0].somModel.tcam_mask[5][624][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][625][0]=80'h00000000db56c981ece6;
sos_loop[0].somModel.tcam_mask[5][625][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][626][0]=80'h00000000cfe8af38f522;
sos_loop[0].somModel.tcam_mask[5][626][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][627][0]=80'h000000008e919d8a745b;
sos_loop[0].somModel.tcam_mask[5][627][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][628][0]=80'h00000000543818958c78;
sos_loop[0].somModel.tcam_mask[5][628][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][629][0]=80'h00000000a8b931f97188;
sos_loop[0].somModel.tcam_mask[5][629][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][630][0]=80'h000000007dee0d849922;
sos_loop[0].somModel.tcam_mask[5][630][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][631][0]=80'h000000001017ca8a2953;
sos_loop[0].somModel.tcam_mask[5][631][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][632][0]=80'h000000007ed9cae24403;
sos_loop[0].somModel.tcam_mask[5][632][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][633][0]=80'h00000000ea187ed4d55a;
sos_loop[0].somModel.tcam_mask[5][633][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][634][0]=80'h000000002e76e28270f1;
sos_loop[0].somModel.tcam_mask[5][634][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][635][0]=80'h00000000f1980343333f;
sos_loop[0].somModel.tcam_mask[5][635][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][636][0]=80'h000000008de1c963c062;
sos_loop[0].somModel.tcam_mask[5][636][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][637][0]=80'h000000003fd86ea44501;
sos_loop[0].somModel.tcam_mask[5][637][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][638][0]=80'h00000000dc791a00bf2c;
sos_loop[0].somModel.tcam_mask[5][638][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][639][0]=80'h0000000076fd772b3105;
sos_loop[0].somModel.tcam_mask[5][639][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][640][0]=80'h000000009137a6d429b2;
sos_loop[0].somModel.tcam_mask[5][640][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][641][0]=80'h0000000049d4cbef7ccc;
sos_loop[0].somModel.tcam_mask[5][641][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][642][0]=80'h000000008051f12b529f;
sos_loop[0].somModel.tcam_mask[5][642][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][643][0]=80'h0000000008d6aa657a5e;
sos_loop[0].somModel.tcam_mask[5][643][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][644][0]=80'h0000000044bafb829ee6;
sos_loop[0].somModel.tcam_mask[5][644][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][645][0]=80'h00000000e55061ccc7b7;
sos_loop[0].somModel.tcam_mask[5][645][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][646][0]=80'h00000000d75970bd3bb0;
sos_loop[0].somModel.tcam_mask[5][646][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][647][0]=80'h000000004811729ba385;
sos_loop[0].somModel.tcam_mask[5][647][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][648][0]=80'h00000000c0501fd955df;
sos_loop[0].somModel.tcam_mask[5][648][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][649][0]=80'h00000000659c29b06d69;
sos_loop[0].somModel.tcam_mask[5][649][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][650][0]=80'h000000006aec373261a3;
sos_loop[0].somModel.tcam_mask[5][650][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][651][0]=80'h00000000c25cd90f5dab;
sos_loop[0].somModel.tcam_mask[5][651][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][652][0]=80'h00000000cee3230bfef6;
sos_loop[0].somModel.tcam_mask[5][652][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][653][0]=80'h000000007bde198a992f;
sos_loop[0].somModel.tcam_mask[5][653][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][654][0]=80'h000000007cd4d9587ccb;
sos_loop[0].somModel.tcam_mask[5][654][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][655][0]=80'h000000005cee7e94dd42;
sos_loop[0].somModel.tcam_mask[5][655][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][656][0]=80'h000000000c7f2c96b613;
sos_loop[0].somModel.tcam_mask[5][656][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][657][0]=80'h00000000f2de9d0bdde4;
sos_loop[0].somModel.tcam_mask[5][657][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][658][0]=80'h00000000b80342294761;
sos_loop[0].somModel.tcam_mask[5][658][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][659][0]=80'h00000000ef05f9051dde;
sos_loop[0].somModel.tcam_mask[5][659][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][660][0]=80'h00000000089d9864b0f7;
sos_loop[0].somModel.tcam_mask[5][660][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[5][661][0]=80'h00000000f84ebc6b5933;
sos_loop[0].somModel.tcam_mask[5][661][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][662][0]=80'h0000000099c7ebd6ef11;
sos_loop[0].somModel.tcam_mask[5][662][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][663][0]=80'h00000000a5cfc726453c;
sos_loop[0].somModel.tcam_mask[5][663][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][664][0]=80'h000000008e33ccc43905;
sos_loop[0].somModel.tcam_mask[5][664][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][665][0]=80'h0000000061dbc393f8b8;
sos_loop[0].somModel.tcam_mask[5][665][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][666][0]=80'h00000000b5776eb8e40c;
sos_loop[0].somModel.tcam_mask[5][666][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][667][0]=80'h00000000c56f02fbb8af;
sos_loop[0].somModel.tcam_mask[5][667][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][668][0]=80'h00000000f06ac89a6e2e;
sos_loop[0].somModel.tcam_mask[5][668][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][669][0]=80'h000000004d46ea5704c7;
sos_loop[0].somModel.tcam_mask[5][669][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][670][0]=80'h00000000018a0d2ab536;
sos_loop[0].somModel.tcam_mask[5][670][0]=80'hfffffffffe0000000000;
sos_loop[0].somModel.tcam_data[5][671][0]=80'h00000000de24ea9c8559;
sos_loop[0].somModel.tcam_mask[5][671][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][672][0]=80'h00000000117c2dcb8a3f;
sos_loop[0].somModel.tcam_mask[5][672][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][673][0]=80'h00000000042c5800a198;
sos_loop[0].somModel.tcam_mask[5][673][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][674][0]=80'h00000000c866641162c8;
sos_loop[0].somModel.tcam_mask[5][674][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][675][0]=80'h00000000c59ce2a178ef;
sos_loop[0].somModel.tcam_mask[5][675][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][676][0]=80'h0000000091b9a88b2186;
sos_loop[0].somModel.tcam_mask[5][676][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][677][0]=80'h00000000baaaa92f9330;
sos_loop[0].somModel.tcam_mask[5][677][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][678][0]=80'h00000000899bc4d45fed;
sos_loop[0].somModel.tcam_mask[5][678][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][679][0]=80'h0000000031aba86c07cd;
sos_loop[0].somModel.tcam_mask[5][679][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][680][0]=80'h00000000c4984e56b9a3;
sos_loop[0].somModel.tcam_mask[5][680][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][681][0]=80'h000000001b2cb5378bd2;
sos_loop[0].somModel.tcam_mask[5][681][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[5][682][0]=80'h00000000ff120ca68f9a;
sos_loop[0].somModel.tcam_mask[5][682][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][683][0]=80'h00000000a835dfd4a64e;
sos_loop[0].somModel.tcam_mask[5][683][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][684][0]=80'h00000000cc35683c57dc;
sos_loop[0].somModel.tcam_mask[5][684][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][685][0]=80'h00000000a5c1099a0ccc;
sos_loop[0].somModel.tcam_mask[5][685][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][686][0]=80'h00000000efd95c4e5fe9;
sos_loop[0].somModel.tcam_mask[5][686][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][687][0]=80'h000000007c76d25796aa;
sos_loop[0].somModel.tcam_mask[5][687][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][688][0]=80'h0000000007b60730923d;
sos_loop[0].somModel.tcam_mask[5][688][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][689][0]=80'h0000000007373b8b8f3c;
sos_loop[0].somModel.tcam_mask[5][689][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[5][690][0]=80'h0000000037e56c799b77;
sos_loop[0].somModel.tcam_mask[5][690][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[5][691][0]=80'h0000000064aeec7ab84c;
sos_loop[0].somModel.tcam_mask[5][691][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][692][0]=80'h00000000dc1814387312;
sos_loop[0].somModel.tcam_mask[5][692][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][693][0]=80'h00000000dd2835b8c4f9;
sos_loop[0].somModel.tcam_mask[5][693][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][694][0]=80'h000000005af2eb552cca;
sos_loop[0].somModel.tcam_mask[5][694][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][695][0]=80'h00000000446b9299fa74;
sos_loop[0].somModel.tcam_mask[5][695][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][696][0]=80'h0000000086928cf64fc6;
sos_loop[0].somModel.tcam_mask[5][696][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][697][0]=80'h00000000c4fdc019c61f;
sos_loop[0].somModel.tcam_mask[5][697][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][698][0]=80'h00000000882f97bb161f;
sos_loop[0].somModel.tcam_mask[5][698][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[5][699][0]=80'h000000004ed606f4518d;
sos_loop[0].somModel.tcam_mask[5][699][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[5][700][0]=80'h00000000bd46a3aa3c15;
sos_loop[0].somModel.tcam_mask[5][700][0]=80'hffffffff000000000000;
sos_loop[0].somModel.sram_dat[5][0][0]=96'hdeadbf;
sos_loop[0].somModel.sram_ptr[5][0]=939;
sos_loop[0].somModel.sram_dat[5][1][0]=96'hec67;
sos_loop[0].somModel.sram_ptr[5][1]=3;
sos_loop[0].somModel.sram_dat[5][2][0]=96'hca33;
sos_loop[0].somModel.sram_ptr[5][2]=3;
sos_loop[0].somModel.sram_dat[5][3][0]=96'h6d67;
sos_loop[0].somModel.sram_ptr[5][3]=3;
sos_loop[0].somModel.sram_dat[5][4][0]=96'hc411;
sos_loop[0].somModel.sram_ptr[5][4]=3;
sos_loop[0].somModel.sram_dat[5][5][0]=96'he871;
sos_loop[0].somModel.sram_ptr[5][5]=3;
sos_loop[0].somModel.sram_dat[5][6][0]=96'h434d;
sos_loop[0].somModel.sram_ptr[5][6]=3;
sos_loop[0].somModel.sram_dat[5][7][0]=96'hbc90;
sos_loop[0].somModel.sram_ptr[5][7]=3;
sos_loop[0].somModel.sram_dat[5][8][0]=96'h3182;
sos_loop[0].somModel.sram_ptr[5][8]=3;
sos_loop[0].somModel.sram_dat[5][9][0]=96'hf995;
sos_loop[0].somModel.sram_ptr[5][9]=3;
sos_loop[0].somModel.sram_dat[5][10][0]=96'hab9b;
sos_loop[0].somModel.sram_ptr[5][10]=3;
sos_loop[0].somModel.sram_dat[5][11][0]=96'h3f0e;
sos_loop[0].somModel.sram_ptr[5][11]=3;
sos_loop[0].somModel.sram_dat[5][12][0]=96'ha49;
sos_loop[0].somModel.sram_ptr[5][12]=3;
sos_loop[0].somModel.sram_dat[5][13][0]=96'h9ced;
sos_loop[0].somModel.sram_ptr[5][13]=3;
sos_loop[0].somModel.sram_dat[5][14][0]=96'hfa16;
sos_loop[0].somModel.sram_ptr[5][14]=3;
sos_loop[0].somModel.sram_dat[5][15][0]=96'hbf3;
sos_loop[0].somModel.sram_ptr[5][15]=3;
sos_loop[0].somModel.sram_dat[5][16][0]=96'hecf9;
sos_loop[0].somModel.sram_ptr[5][16]=3;
sos_loop[0].somModel.sram_dat[5][17][0]=96'h273b;
sos_loop[0].somModel.sram_ptr[5][17]=3;
sos_loop[0].somModel.sram_dat[5][18][0]=96'h7d62;
sos_loop[0].somModel.sram_ptr[5][18]=3;
sos_loop[0].somModel.sram_dat[5][19][0]=96'h3658;
sos_loop[0].somModel.sram_ptr[5][19]=3;
sos_loop[0].somModel.sram_dat[5][20][0]=96'hd34c;
sos_loop[0].somModel.sram_ptr[5][20]=3;
sos_loop[0].somModel.sram_dat[5][21][0]=96'ha11e;
sos_loop[0].somModel.sram_ptr[5][21]=3;
sos_loop[0].somModel.sram_dat[5][22][0]=96'hcdb1;
sos_loop[0].somModel.sram_ptr[5][22]=3;
sos_loop[0].somModel.sram_dat[5][23][0]=96'hcb23;
sos_loop[0].somModel.sram_ptr[5][23]=3;
sos_loop[0].somModel.sram_dat[5][24][0]=96'h4f15;
sos_loop[0].somModel.sram_ptr[5][24]=3;
sos_loop[0].somModel.sram_dat[5][25][0]=96'hf6;
sos_loop[0].somModel.sram_ptr[5][25]=3;
sos_loop[0].somModel.sram_dat[5][26][0]=96'h8a2b;
sos_loop[0].somModel.sram_ptr[5][26]=3;
sos_loop[0].somModel.sram_dat[5][27][0]=96'hb21;
sos_loop[0].somModel.sram_ptr[5][27]=3;
sos_loop[0].somModel.sram_dat[5][28][0]=96'h1699;
sos_loop[0].somModel.sram_ptr[5][28]=3;
sos_loop[0].somModel.sram_dat[5][29][0]=96'h1d0;
sos_loop[0].somModel.sram_ptr[5][29]=3;
sos_loop[0].somModel.sram_dat[5][30][0]=96'hdaf2;
sos_loop[0].somModel.sram_ptr[5][30]=3;
sos_loop[0].somModel.sram_dat[5][31][0]=96'h317c;
sos_loop[0].somModel.sram_ptr[5][31]=3;
sos_loop[0].somModel.sram_dat[5][32][0]=96'h5312;
sos_loop[0].somModel.sram_ptr[5][32]=3;
sos_loop[0].somModel.sram_dat[5][33][0]=96'hcd1a;
sos_loop[0].somModel.sram_ptr[5][33]=3;
sos_loop[0].somModel.sram_dat[5][34][0]=96'h24e6;
sos_loop[0].somModel.sram_ptr[5][34]=3;
sos_loop[0].somModel.sram_dat[5][35][0]=96'h8650;
sos_loop[0].somModel.sram_ptr[5][35]=3;
sos_loop[0].somModel.sram_dat[5][36][0]=96'h948a;
sos_loop[0].somModel.sram_ptr[5][36]=3;
sos_loop[0].somModel.sram_dat[5][37][0]=96'h3b16;
sos_loop[0].somModel.sram_ptr[5][37]=3;
sos_loop[0].somModel.sram_dat[5][38][0]=96'hd1cc;
sos_loop[0].somModel.sram_ptr[5][38]=3;
sos_loop[0].somModel.sram_dat[5][39][0]=96'hed39;
sos_loop[0].somModel.sram_ptr[5][39]=3;
sos_loop[0].somModel.sram_dat[5][40][0]=96'h4552;
sos_loop[0].somModel.sram_ptr[5][40]=3;
sos_loop[0].somModel.sram_dat[5][41][0]=96'h3604;
sos_loop[0].somModel.sram_ptr[5][41]=3;
sos_loop[0].somModel.sram_dat[5][42][0]=96'h128b;
sos_loop[0].somModel.sram_ptr[5][42]=3;
sos_loop[0].somModel.sram_dat[5][43][0]=96'he052;
sos_loop[0].somModel.sram_ptr[5][43]=3;
sos_loop[0].somModel.sram_dat[5][44][0]=96'h9626;
sos_loop[0].somModel.sram_ptr[5][44]=3;
sos_loop[0].somModel.sram_dat[5][45][0]=96'h6ae6;
sos_loop[0].somModel.sram_ptr[5][45]=3;
sos_loop[0].somModel.sram_dat[5][46][0]=96'h5c87;
sos_loop[0].somModel.sram_ptr[5][46]=3;
sos_loop[0].somModel.sram_dat[5][47][0]=96'h8b78;
sos_loop[0].somModel.sram_ptr[5][47]=3;
sos_loop[0].somModel.sram_dat[5][48][0]=96'h4875;
sos_loop[0].somModel.sram_ptr[5][48]=3;
sos_loop[0].somModel.sram_dat[5][49][0]=96'h2d1e;
sos_loop[0].somModel.sram_ptr[5][49]=3;
sos_loop[0].somModel.sram_dat[5][50][0]=96'h5b49;
sos_loop[0].somModel.sram_ptr[5][50]=3;
sos_loop[0].somModel.sram_dat[5][51][0]=96'h59b7;
sos_loop[0].somModel.sram_ptr[5][51]=3;
sos_loop[0].somModel.sram_dat[5][52][0]=96'he851;
sos_loop[0].somModel.sram_ptr[5][52]=3;
sos_loop[0].somModel.sram_dat[5][53][0]=96'h5ca1;
sos_loop[0].somModel.sram_ptr[5][53]=3;
sos_loop[0].somModel.sram_dat[5][54][0]=96'h7ba3;
sos_loop[0].somModel.sram_ptr[5][54]=3;
sos_loop[0].somModel.sram_dat[5][55][0]=96'h2c4;
sos_loop[0].somModel.sram_ptr[5][55]=3;
sos_loop[0].somModel.sram_dat[5][56][0]=96'h4df4;
sos_loop[0].somModel.sram_ptr[5][56]=3;
sos_loop[0].somModel.sram_dat[5][57][0]=96'h6933;
sos_loop[0].somModel.sram_ptr[5][57]=3;
sos_loop[0].somModel.sram_dat[5][58][0]=96'he4f4;
sos_loop[0].somModel.sram_ptr[5][58]=3;
sos_loop[0].somModel.sram_dat[5][59][0]=96'he474;
sos_loop[0].somModel.sram_ptr[5][59]=3;
sos_loop[0].somModel.sram_dat[5][60][0]=96'hb8d7;
sos_loop[0].somModel.sram_ptr[5][60]=3;
sos_loop[0].somModel.sram_dat[5][61][0]=96'h3227;
sos_loop[0].somModel.sram_ptr[5][61]=3;
sos_loop[0].somModel.sram_dat[5][62][0]=96'haae6;
sos_loop[0].somModel.sram_ptr[5][62]=3;
sos_loop[0].somModel.sram_dat[5][63][0]=96'h62c4;
sos_loop[0].somModel.sram_ptr[5][63]=3;
sos_loop[0].somModel.sram_dat[5][64][0]=96'hdd68;
sos_loop[0].somModel.sram_ptr[5][64]=3;
sos_loop[0].somModel.sram_dat[5][65][0]=96'h7e73;
sos_loop[0].somModel.sram_ptr[5][65]=3;
sos_loop[0].somModel.sram_dat[5][66][0]=96'h3af;
sos_loop[0].somModel.sram_ptr[5][66]=3;
sos_loop[0].somModel.sram_dat[5][67][0]=96'h48de;
sos_loop[0].somModel.sram_ptr[5][67]=3;
sos_loop[0].somModel.sram_dat[5][68][0]=96'hefd;
sos_loop[0].somModel.sram_ptr[5][68]=3;
sos_loop[0].somModel.sram_dat[5][69][0]=96'he419;
sos_loop[0].somModel.sram_ptr[5][69]=3;
sos_loop[0].somModel.sram_dat[5][70][0]=96'h9356;
sos_loop[0].somModel.sram_ptr[5][70]=3;
sos_loop[0].somModel.sram_dat[5][71][0]=96'ha8b9;
sos_loop[0].somModel.sram_ptr[5][71]=3;
sos_loop[0].somModel.sram_dat[5][72][0]=96'h64c1;
sos_loop[0].somModel.sram_ptr[5][72]=3;
sos_loop[0].somModel.sram_dat[5][73][0]=96'hb6da;
sos_loop[0].somModel.sram_ptr[5][73]=3;
sos_loop[0].somModel.sram_dat[5][74][0]=96'hea32;
sos_loop[0].somModel.sram_ptr[5][74]=3;
sos_loop[0].somModel.sram_dat[5][75][0]=96'h5eed;
sos_loop[0].somModel.sram_ptr[5][75]=3;
sos_loop[0].somModel.sram_dat[5][76][0]=96'hfaf4;
sos_loop[0].somModel.sram_ptr[5][76]=3;
sos_loop[0].somModel.sram_dat[5][77][0]=96'h7a2c;
sos_loop[0].somModel.sram_ptr[5][77]=3;
sos_loop[0].somModel.sram_dat[5][78][0]=96'hf957;
sos_loop[0].somModel.sram_ptr[5][78]=3;
sos_loop[0].somModel.sram_dat[5][79][0]=96'h5b6b;
sos_loop[0].somModel.sram_ptr[5][79]=3;
sos_loop[0].somModel.sram_dat[5][80][0]=96'h3d98;
sos_loop[0].somModel.sram_ptr[5][80]=3;
sos_loop[0].somModel.sram_dat[5][81][0]=96'hf6bf;
sos_loop[0].somModel.sram_ptr[5][81]=3;
sos_loop[0].somModel.sram_dat[5][82][0]=96'h933e;
sos_loop[0].somModel.sram_ptr[5][82]=3;
sos_loop[0].somModel.sram_dat[5][83][0]=96'h4e1f;
sos_loop[0].somModel.sram_ptr[5][83]=3;
sos_loop[0].somModel.sram_dat[5][84][0]=96'h7a3d;
sos_loop[0].somModel.sram_ptr[5][84]=3;
sos_loop[0].somModel.sram_dat[5][85][0]=96'h7d64;
sos_loop[0].somModel.sram_ptr[5][85]=3;
sos_loop[0].somModel.sram_dat[5][86][0]=96'hdfa6;
sos_loop[0].somModel.sram_ptr[5][86]=3;
sos_loop[0].somModel.sram_dat[5][87][0]=96'he19a;
sos_loop[0].somModel.sram_ptr[5][87]=3;
sos_loop[0].somModel.sram_dat[5][88][0]=96'h66d1;
sos_loop[0].somModel.sram_ptr[5][88]=3;
sos_loop[0].somModel.sram_dat[5][89][0]=96'hf6c4;
sos_loop[0].somModel.sram_ptr[5][89]=3;
sos_loop[0].somModel.sram_dat[5][90][0]=96'hacc9;
sos_loop[0].somModel.sram_ptr[5][90]=3;
sos_loop[0].somModel.sram_dat[5][91][0]=96'ha5aa;
sos_loop[0].somModel.sram_ptr[5][91]=3;
sos_loop[0].somModel.sram_dat[5][92][0]=96'h777f;
sos_loop[0].somModel.sram_ptr[5][92]=3;
sos_loop[0].somModel.sram_dat[5][93][0]=96'hf0f0;
sos_loop[0].somModel.sram_ptr[5][93]=3;
sos_loop[0].somModel.sram_dat[5][94][0]=96'hcfbb;
sos_loop[0].somModel.sram_ptr[5][94]=3;
sos_loop[0].somModel.sram_dat[5][95][0]=96'h2c19;
sos_loop[0].somModel.sram_ptr[5][95]=3;
sos_loop[0].somModel.sram_dat[5][96][0]=96'h24d4;
sos_loop[0].somModel.sram_ptr[5][96]=3;
sos_loop[0].somModel.sram_dat[5][97][0]=96'h5ffc;
sos_loop[0].somModel.sram_ptr[5][97]=3;
sos_loop[0].somModel.sram_dat[5][98][0]=96'hacf5;
sos_loop[0].somModel.sram_ptr[5][98]=3;
sos_loop[0].somModel.sram_dat[5][99][0]=96'h894c;
sos_loop[0].somModel.sram_ptr[5][99]=3;
sos_loop[0].somModel.sram_dat[5][100][0]=96'h17ab;
sos_loop[0].somModel.sram_ptr[5][100]=3;
sos_loop[0].somModel.sram_dat[5][101][0]=96'h1075;
sos_loop[0].somModel.sram_ptr[5][101]=3;
sos_loop[0].somModel.sram_dat[5][102][0]=96'h5677;
sos_loop[0].somModel.sram_ptr[5][102]=3;
sos_loop[0].somModel.sram_dat[5][103][0]=96'h1b39;
sos_loop[0].somModel.sram_ptr[5][103]=3;
sos_loop[0].somModel.sram_dat[5][104][0]=96'h3a80;
sos_loop[0].somModel.sram_ptr[5][104]=3;
sos_loop[0].somModel.sram_dat[5][105][0]=96'h3017;
sos_loop[0].somModel.sram_ptr[5][105]=3;
sos_loop[0].somModel.sram_dat[5][106][0]=96'h9202;
sos_loop[0].somModel.sram_ptr[5][106]=3;
sos_loop[0].somModel.sram_dat[5][107][0]=96'h74cd;
sos_loop[0].somModel.sram_ptr[5][107]=3;
sos_loop[0].somModel.sram_dat[5][108][0]=96'h5c5f;
sos_loop[0].somModel.sram_ptr[5][108]=3;
sos_loop[0].somModel.sram_dat[5][109][0]=96'h1117;
sos_loop[0].somModel.sram_ptr[5][109]=3;
sos_loop[0].somModel.sram_dat[5][110][0]=96'he794;
sos_loop[0].somModel.sram_ptr[5][110]=3;
sos_loop[0].somModel.sram_dat[5][111][0]=96'ha456;
sos_loop[0].somModel.sram_ptr[5][111]=3;
sos_loop[0].somModel.sram_dat[5][112][0]=96'hcfdd;
sos_loop[0].somModel.sram_ptr[5][112]=3;
sos_loop[0].somModel.sram_dat[5][113][0]=96'hd835;
sos_loop[0].somModel.sram_ptr[5][113]=3;
sos_loop[0].somModel.sram_dat[5][114][0]=96'hdd49;
sos_loop[0].somModel.sram_ptr[5][114]=3;
sos_loop[0].somModel.sram_dat[5][115][0]=96'h7570;
sos_loop[0].somModel.sram_ptr[5][115]=3;
sos_loop[0].somModel.sram_dat[5][116][0]=96'hb255;
sos_loop[0].somModel.sram_ptr[5][116]=3;
sos_loop[0].somModel.sram_dat[5][117][0]=96'h6980;
sos_loop[0].somModel.sram_ptr[5][117]=3;
sos_loop[0].somModel.sram_dat[5][118][0]=96'h8260;
sos_loop[0].somModel.sram_ptr[5][118]=3;
sos_loop[0].somModel.sram_dat[5][119][0]=96'ha205;
sos_loop[0].somModel.sram_ptr[5][119]=3;
sos_loop[0].somModel.sram_dat[5][120][0]=96'h304d;
sos_loop[0].somModel.sram_ptr[5][120]=3;
sos_loop[0].somModel.sram_dat[5][121][0]=96'hfb08;
sos_loop[0].somModel.sram_ptr[5][121]=3;
sos_loop[0].somModel.sram_dat[5][122][0]=96'hfa71;
sos_loop[0].somModel.sram_ptr[5][122]=3;
sos_loop[0].somModel.sram_dat[5][123][0]=96'he4d8;
sos_loop[0].somModel.sram_ptr[5][123]=3;
sos_loop[0].somModel.sram_dat[5][124][0]=96'h1c3e;
sos_loop[0].somModel.sram_ptr[5][124]=3;
sos_loop[0].somModel.sram_dat[5][125][0]=96'h4931;
sos_loop[0].somModel.sram_ptr[5][125]=3;
sos_loop[0].somModel.sram_dat[5][126][0]=96'h84b5;
sos_loop[0].somModel.sram_ptr[5][126]=3;
sos_loop[0].somModel.sram_dat[5][127][0]=96'h711;
sos_loop[0].somModel.sram_ptr[5][127]=3;
sos_loop[0].somModel.sram_dat[5][128][0]=96'hca64;
sos_loop[0].somModel.sram_ptr[5][128]=3;
sos_loop[0].somModel.sram_dat[5][129][0]=96'hd669;
sos_loop[0].somModel.sram_ptr[5][129]=3;
sos_loop[0].somModel.sram_dat[5][130][0]=96'h4363;
sos_loop[0].somModel.sram_ptr[5][130]=3;
sos_loop[0].somModel.sram_dat[5][131][0]=96'hf838;
sos_loop[0].somModel.sram_ptr[5][131]=3;
sos_loop[0].somModel.sram_dat[5][132][0]=96'h8a28;
sos_loop[0].somModel.sram_ptr[5][132]=3;
sos_loop[0].somModel.sram_dat[5][133][0]=96'h811a;
sos_loop[0].somModel.sram_ptr[5][133]=3;
sos_loop[0].somModel.sram_dat[5][134][0]=96'h40c;
sos_loop[0].somModel.sram_ptr[5][134]=3;
sos_loop[0].somModel.sram_dat[5][135][0]=96'h41ac;
sos_loop[0].somModel.sram_ptr[5][135]=3;
sos_loop[0].somModel.sram_dat[5][136][0]=96'h4b1b;
sos_loop[0].somModel.sram_ptr[5][136]=3;
sos_loop[0].somModel.sram_dat[5][137][0]=96'hb214;
sos_loop[0].somModel.sram_ptr[5][137]=3;
sos_loop[0].somModel.sram_dat[5][138][0]=96'h504f;
sos_loop[0].somModel.sram_ptr[5][138]=3;
sos_loop[0].somModel.sram_dat[5][139][0]=96'hae5d;
sos_loop[0].somModel.sram_ptr[5][139]=3;
sos_loop[0].somModel.sram_dat[5][140][0]=96'h914b;
sos_loop[0].somModel.sram_ptr[5][140]=3;
sos_loop[0].somModel.sram_dat[5][141][0]=96'h4c67;
sos_loop[0].somModel.sram_ptr[5][141]=3;
sos_loop[0].somModel.sram_dat[5][142][0]=96'h25f9;
sos_loop[0].somModel.sram_ptr[5][142]=3;
sos_loop[0].somModel.sram_dat[5][143][0]=96'h2323;
sos_loop[0].somModel.sram_ptr[5][143]=3;
sos_loop[0].somModel.sram_dat[5][144][0]=96'h3f89;
sos_loop[0].somModel.sram_ptr[5][144]=3;
sos_loop[0].somModel.sram_dat[5][145][0]=96'h5c3;
sos_loop[0].somModel.sram_ptr[5][145]=3;
sos_loop[0].somModel.sram_dat[5][146][0]=96'h8362;
sos_loop[0].somModel.sram_ptr[5][146]=3;
sos_loop[0].somModel.sram_dat[5][147][0]=96'hd4ed;
sos_loop[0].somModel.sram_ptr[5][147]=3;
sos_loop[0].somModel.sram_dat[5][148][0]=96'h1634;
sos_loop[0].somModel.sram_ptr[5][148]=3;
sos_loop[0].somModel.sram_dat[5][149][0]=96'h6bb4;
sos_loop[0].somModel.sram_ptr[5][149]=3;
sos_loop[0].somModel.sram_dat[5][150][0]=96'h8ca3;
sos_loop[0].somModel.sram_ptr[5][150]=3;
sos_loop[0].somModel.sram_dat[5][151][0]=96'hc978;
sos_loop[0].somModel.sram_ptr[5][151]=3;
sos_loop[0].somModel.sram_dat[5][152][0]=96'hf216;
sos_loop[0].somModel.sram_ptr[5][152]=3;
sos_loop[0].somModel.sram_dat[5][153][0]=96'hcd29;
sos_loop[0].somModel.sram_ptr[5][153]=3;
sos_loop[0].somModel.sram_dat[5][154][0]=96'h5114;
sos_loop[0].somModel.sram_ptr[5][154]=3;
sos_loop[0].somModel.sram_dat[5][155][0]=96'h5ffc;
sos_loop[0].somModel.sram_ptr[5][155]=3;
sos_loop[0].somModel.sram_dat[5][156][0]=96'hefa8;
sos_loop[0].somModel.sram_ptr[5][156]=3;
sos_loop[0].somModel.sram_dat[5][157][0]=96'ha3;
sos_loop[0].somModel.sram_ptr[5][157]=3;
sos_loop[0].somModel.sram_dat[5][158][0]=96'h5bcb;
sos_loop[0].somModel.sram_ptr[5][158]=3;
sos_loop[0].somModel.sram_dat[5][159][0]=96'h34d2;
sos_loop[0].somModel.sram_ptr[5][159]=3;
sos_loop[0].somModel.sram_dat[5][160][0]=96'hb6ed;
sos_loop[0].somModel.sram_ptr[5][160]=3;
sos_loop[0].somModel.sram_dat[5][161][0]=96'h2d7a;
sos_loop[0].somModel.sram_ptr[5][161]=3;
sos_loop[0].somModel.sram_dat[5][162][0]=96'h53b8;
sos_loop[0].somModel.sram_ptr[5][162]=3;
sos_loop[0].somModel.sram_dat[5][163][0]=96'h9151;
sos_loop[0].somModel.sram_ptr[5][163]=3;
sos_loop[0].somModel.sram_dat[5][164][0]=96'h8bc6;
sos_loop[0].somModel.sram_ptr[5][164]=3;
sos_loop[0].somModel.sram_dat[5][165][0]=96'h74ce;
sos_loop[0].somModel.sram_ptr[5][165]=3;
sos_loop[0].somModel.sram_dat[5][166][0]=96'h300e;
sos_loop[0].somModel.sram_ptr[5][166]=3;
sos_loop[0].somModel.sram_dat[5][167][0]=96'h6347;
sos_loop[0].somModel.sram_ptr[5][167]=3;
sos_loop[0].somModel.sram_dat[5][168][0]=96'h8a2f;
sos_loop[0].somModel.sram_ptr[5][168]=3;
sos_loop[0].somModel.sram_dat[5][169][0]=96'h775b;
sos_loop[0].somModel.sram_ptr[5][169]=3;
sos_loop[0].somModel.sram_dat[5][170][0]=96'hb202;
sos_loop[0].somModel.sram_ptr[5][170]=3;
sos_loop[0].somModel.sram_dat[5][171][0]=96'h43c7;
sos_loop[0].somModel.sram_ptr[5][171]=3;
sos_loop[0].somModel.sram_dat[5][172][0]=96'h77bb;
sos_loop[0].somModel.sram_ptr[5][172]=3;
sos_loop[0].somModel.sram_dat[5][173][0]=96'h567e;
sos_loop[0].somModel.sram_ptr[5][173]=3;
sos_loop[0].somModel.sram_dat[5][174][0]=96'h8d37;
sos_loop[0].somModel.sram_ptr[5][174]=3;
sos_loop[0].somModel.sram_dat[5][175][0]=96'hf369;
sos_loop[0].somModel.sram_ptr[5][175]=3;
sos_loop[0].somModel.sram_dat[5][176][0]=96'h3a0f;
sos_loop[0].somModel.sram_ptr[5][176]=3;
sos_loop[0].somModel.sram_dat[5][177][0]=96'ha1f5;
sos_loop[0].somModel.sram_ptr[5][177]=3;
sos_loop[0].somModel.sram_dat[5][178][0]=96'h76a9;
sos_loop[0].somModel.sram_ptr[5][178]=3;
sos_loop[0].somModel.sram_dat[5][179][0]=96'h1474;
sos_loop[0].somModel.sram_ptr[5][179]=3;
sos_loop[0].somModel.sram_dat[5][180][0]=96'h52e6;
sos_loop[0].somModel.sram_ptr[5][180]=3;
sos_loop[0].somModel.sram_dat[5][181][0]=96'h2f51;
sos_loop[0].somModel.sram_ptr[5][181]=3;
sos_loop[0].somModel.sram_dat[5][182][0]=96'h652b;
sos_loop[0].somModel.sram_ptr[5][182]=3;
sos_loop[0].somModel.sram_dat[5][183][0]=96'he3f9;
sos_loop[0].somModel.sram_ptr[5][183]=3;
sos_loop[0].somModel.sram_dat[5][184][0]=96'ha7a;
sos_loop[0].somModel.sram_ptr[5][184]=3;
sos_loop[0].somModel.sram_dat[5][185][0]=96'hb249;
sos_loop[0].somModel.sram_ptr[5][185]=3;
sos_loop[0].somModel.sram_dat[5][186][0]=96'h32a0;
sos_loop[0].somModel.sram_ptr[5][186]=3;
sos_loop[0].somModel.sram_dat[5][187][0]=96'h6074;
sos_loop[0].somModel.sram_ptr[5][187]=3;
sos_loop[0].somModel.sram_dat[5][188][0]=96'h3737;
sos_loop[0].somModel.sram_ptr[5][188]=3;
sos_loop[0].somModel.sram_dat[5][189][0]=96'h2dfa;
sos_loop[0].somModel.sram_ptr[5][189]=3;
sos_loop[0].somModel.sram_dat[5][190][0]=96'ha1f2;
sos_loop[0].somModel.sram_ptr[5][190]=3;
sos_loop[0].somModel.sram_dat[5][191][0]=96'h4653;
sos_loop[0].somModel.sram_ptr[5][191]=3;
sos_loop[0].somModel.sram_dat[5][192][0]=96'h27fb;
sos_loop[0].somModel.sram_ptr[5][192]=3;
sos_loop[0].somModel.sram_dat[5][193][0]=96'he2cf;
sos_loop[0].somModel.sram_ptr[5][193]=3;
sos_loop[0].somModel.sram_dat[5][194][0]=96'hc65c;
sos_loop[0].somModel.sram_ptr[5][194]=3;
sos_loop[0].somModel.sram_dat[5][195][0]=96'hcfb9;
sos_loop[0].somModel.sram_ptr[5][195]=3;
sos_loop[0].somModel.sram_dat[5][196][0]=96'h295;
sos_loop[0].somModel.sram_ptr[5][196]=3;
sos_loop[0].somModel.sram_dat[5][197][0]=96'h639d;
sos_loop[0].somModel.sram_ptr[5][197]=3;
sos_loop[0].somModel.sram_dat[5][198][0]=96'h7807;
sos_loop[0].somModel.sram_ptr[5][198]=3;
sos_loop[0].somModel.sram_dat[5][199][0]=96'h14ab;
sos_loop[0].somModel.sram_ptr[5][199]=3;
sos_loop[0].somModel.sram_dat[5][200][0]=96'h2540;
sos_loop[0].somModel.sram_ptr[5][200]=3;
sos_loop[0].somModel.sram_dat[5][201][0]=96'ha6b5;
sos_loop[0].somModel.sram_ptr[5][201]=3;
sos_loop[0].somModel.sram_dat[5][202][0]=96'h349d;
sos_loop[0].somModel.sram_ptr[5][202]=3;
sos_loop[0].somModel.sram_dat[5][203][0]=96'hd281;
sos_loop[0].somModel.sram_ptr[5][203]=3;
sos_loop[0].somModel.sram_dat[5][204][0]=96'h142d;
sos_loop[0].somModel.sram_ptr[5][204]=3;
sos_loop[0].somModel.sram_dat[5][205][0]=96'h6d0d;
sos_loop[0].somModel.sram_ptr[5][205]=3;
sos_loop[0].somModel.sram_dat[5][206][0]=96'he636;
sos_loop[0].somModel.sram_ptr[5][206]=3;
sos_loop[0].somModel.sram_dat[5][207][0]=96'ha342;
sos_loop[0].somModel.sram_ptr[5][207]=3;
sos_loop[0].somModel.sram_dat[5][208][0]=96'h25d3;
sos_loop[0].somModel.sram_ptr[5][208]=3;
sos_loop[0].somModel.sram_dat[5][209][0]=96'hacf;
sos_loop[0].somModel.sram_ptr[5][209]=3;
sos_loop[0].somModel.sram_dat[5][210][0]=96'h58ca;
sos_loop[0].somModel.sram_ptr[5][210]=3;
sos_loop[0].somModel.sram_dat[5][211][0]=96'hb00e;
sos_loop[0].somModel.sram_ptr[5][211]=3;
sos_loop[0].somModel.sram_dat[5][212][0]=96'hb9c1;
sos_loop[0].somModel.sram_ptr[5][212]=3;
sos_loop[0].somModel.sram_dat[5][213][0]=96'h91d;
sos_loop[0].somModel.sram_ptr[5][213]=3;
sos_loop[0].somModel.sram_dat[5][214][0]=96'h8e15;
sos_loop[0].somModel.sram_ptr[5][214]=3;
sos_loop[0].somModel.sram_dat[5][215][0]=96'hff14;
sos_loop[0].somModel.sram_ptr[5][215]=3;
sos_loop[0].somModel.sram_dat[5][216][0]=96'h57fa;
sos_loop[0].somModel.sram_ptr[5][216]=3;
sos_loop[0].somModel.sram_dat[5][217][0]=96'hda3f;
sos_loop[0].somModel.sram_ptr[5][217]=3;
sos_loop[0].somModel.sram_dat[5][218][0]=96'hf47;
sos_loop[0].somModel.sram_ptr[5][218]=3;
sos_loop[0].somModel.sram_dat[5][219][0]=96'had05;
sos_loop[0].somModel.sram_ptr[5][219]=3;
sos_loop[0].somModel.sram_dat[5][220][0]=96'h5563;
sos_loop[0].somModel.sram_ptr[5][220]=3;
sos_loop[0].somModel.sram_dat[5][221][0]=96'h534f;
sos_loop[0].somModel.sram_ptr[5][221]=3;
sos_loop[0].somModel.sram_dat[5][222][0]=96'h327f;
sos_loop[0].somModel.sram_ptr[5][222]=3;
sos_loop[0].somModel.sram_dat[5][223][0]=96'h7e5b;
sos_loop[0].somModel.sram_ptr[5][223]=3;
sos_loop[0].somModel.sram_dat[5][224][0]=96'hadda;
sos_loop[0].somModel.sram_ptr[5][224]=3;
sos_loop[0].somModel.sram_dat[5][225][0]=96'hc981;
sos_loop[0].somModel.sram_ptr[5][225]=3;
sos_loop[0].somModel.sram_dat[5][226][0]=96'hd139;
sos_loop[0].somModel.sram_ptr[5][226]=3;
sos_loop[0].somModel.sram_dat[5][227][0]=96'h2513;
sos_loop[0].somModel.sram_ptr[5][227]=3;
sos_loop[0].somModel.sram_dat[5][228][0]=96'h327d;
sos_loop[0].somModel.sram_ptr[5][228]=3;
sos_loop[0].somModel.sram_dat[5][229][0]=96'h9e05;
sos_loop[0].somModel.sram_ptr[5][229]=3;
sos_loop[0].somModel.sram_dat[5][230][0]=96'hf241;
sos_loop[0].somModel.sram_ptr[5][230]=3;
sos_loop[0].somModel.sram_dat[5][231][0]=96'h1dee;
sos_loop[0].somModel.sram_ptr[5][231]=3;
sos_loop[0].somModel.sram_dat[5][232][0]=96'hd55e;
sos_loop[0].somModel.sram_ptr[5][232]=3;
sos_loop[0].somModel.sram_dat[5][233][0]=96'h25de;
sos_loop[0].somModel.sram_ptr[5][233]=3;
sos_loop[0].somModel.sram_dat[5][234][0]=96'hdf66;
sos_loop[0].somModel.sram_ptr[5][234]=3;
sos_loop[0].somModel.sram_dat[5][235][0]=96'h260e;
sos_loop[0].somModel.sram_ptr[5][235]=3;
sos_loop[0].somModel.sram_dat[5][236][0]=96'h11f9;
sos_loop[0].somModel.sram_ptr[5][236]=3;
sos_loop[0].somModel.sram_dat[5][237][0]=96'h7851;
sos_loop[0].somModel.sram_ptr[5][237]=3;
sos_loop[0].somModel.sram_dat[5][238][0]=96'h4bb5;
sos_loop[0].somModel.sram_ptr[5][238]=3;
sos_loop[0].somModel.sram_dat[5][239][0]=96'h58ad;
sos_loop[0].somModel.sram_ptr[5][239]=3;
sos_loop[0].somModel.sram_dat[5][240][0]=96'hcd39;
sos_loop[0].somModel.sram_ptr[5][240]=3;
sos_loop[0].somModel.sram_dat[5][241][0]=96'h4594;
sos_loop[0].somModel.sram_ptr[5][241]=3;
sos_loop[0].somModel.sram_dat[5][242][0]=96'h9e8b;
sos_loop[0].somModel.sram_ptr[5][242]=3;
sos_loop[0].somModel.sram_dat[5][243][0]=96'h7e25;
sos_loop[0].somModel.sram_ptr[5][243]=3;
sos_loop[0].somModel.sram_dat[5][244][0]=96'h9c66;
sos_loop[0].somModel.sram_ptr[5][244]=3;
sos_loop[0].somModel.sram_dat[5][245][0]=96'h67e;
sos_loop[0].somModel.sram_ptr[5][245]=3;
sos_loop[0].somModel.sram_dat[5][246][0]=96'h1f05;
sos_loop[0].somModel.sram_ptr[5][246]=3;
sos_loop[0].somModel.sram_dat[5][247][0]=96'h3663;
sos_loop[0].somModel.sram_ptr[5][247]=3;
sos_loop[0].somModel.sram_dat[5][248][0]=96'hc3fb;
sos_loop[0].somModel.sram_ptr[5][248]=3;
sos_loop[0].somModel.sram_dat[5][249][0]=96'h689d;
sos_loop[0].somModel.sram_ptr[5][249]=3;
sos_loop[0].somModel.sram_dat[5][250][0]=96'h6519;
sos_loop[0].somModel.sram_ptr[5][250]=3;
sos_loop[0].somModel.sram_dat[5][251][0]=96'hefd8;
sos_loop[0].somModel.sram_ptr[5][251]=3;
sos_loop[0].somModel.sram_dat[5][252][0]=96'hcf65;
sos_loop[0].somModel.sram_ptr[5][252]=3;
sos_loop[0].somModel.sram_dat[5][253][0]=96'h2090;
sos_loop[0].somModel.sram_ptr[5][253]=3;
sos_loop[0].somModel.sram_dat[5][254][0]=96'h7423;
sos_loop[0].somModel.sram_ptr[5][254]=3;
sos_loop[0].somModel.sram_dat[5][255][0]=96'h2ac0;
sos_loop[0].somModel.sram_ptr[5][255]=3;
sos_loop[0].somModel.sram_dat[5][256][0]=96'h5ce1;
sos_loop[0].somModel.sram_ptr[5][256]=3;
sos_loop[0].somModel.sram_dat[5][257][0]=96'h2f49;
sos_loop[0].somModel.sram_ptr[5][257]=3;
sos_loop[0].somModel.sram_dat[5][258][0]=96'he74d;
sos_loop[0].somModel.sram_ptr[5][258]=3;
sos_loop[0].somModel.sram_dat[5][259][0]=96'hfe3a;
sos_loop[0].somModel.sram_ptr[5][259]=3;
sos_loop[0].somModel.sram_dat[5][260][0]=96'h1570;
sos_loop[0].somModel.sram_ptr[5][260]=3;
sos_loop[0].somModel.sram_dat[5][261][0]=96'h96ed;
sos_loop[0].somModel.sram_ptr[5][261]=3;
sos_loop[0].somModel.sram_dat[5][262][0]=96'h2b86;
sos_loop[0].somModel.sram_ptr[5][262]=3;
sos_loop[0].somModel.sram_dat[5][263][0]=96'h3c2;
sos_loop[0].somModel.sram_ptr[5][263]=3;
sos_loop[0].somModel.sram_dat[5][264][0]=96'hd542;
sos_loop[0].somModel.sram_ptr[5][264]=3;
sos_loop[0].somModel.sram_dat[5][265][0]=96'h5df5;
sos_loop[0].somModel.sram_ptr[5][265]=3;
sos_loop[0].somModel.sram_dat[5][266][0]=96'h8aa0;
sos_loop[0].somModel.sram_ptr[5][266]=3;
sos_loop[0].somModel.sram_dat[5][267][0]=96'ha9a3;
sos_loop[0].somModel.sram_ptr[5][267]=3;
sos_loop[0].somModel.sram_dat[5][268][0]=96'h42d3;
sos_loop[0].somModel.sram_ptr[5][268]=3;
sos_loop[0].somModel.sram_dat[5][269][0]=96'h8837;
sos_loop[0].somModel.sram_ptr[5][269]=3;
sos_loop[0].somModel.sram_dat[5][270][0]=96'h3ced;
sos_loop[0].somModel.sram_ptr[5][270]=3;
sos_loop[0].somModel.sram_dat[5][271][0]=96'h48b0;
sos_loop[0].somModel.sram_ptr[5][271]=3;
sos_loop[0].somModel.sram_dat[5][272][0]=96'hd5f;
sos_loop[0].somModel.sram_ptr[5][272]=3;
sos_loop[0].somModel.sram_dat[5][273][0]=96'hf9fd;
sos_loop[0].somModel.sram_ptr[5][273]=3;
sos_loop[0].somModel.sram_dat[5][274][0]=96'h12ac;
sos_loop[0].somModel.sram_ptr[5][274]=3;
sos_loop[0].somModel.sram_dat[5][275][0]=96'h9222;
sos_loop[0].somModel.sram_ptr[5][275]=3;
sos_loop[0].somModel.sram_dat[5][276][0]=96'h4182;
sos_loop[0].somModel.sram_ptr[5][276]=3;
sos_loop[0].somModel.sram_dat[5][277][0]=96'h9201;
sos_loop[0].somModel.sram_ptr[5][277]=3;
sos_loop[0].somModel.sram_dat[5][278][0]=96'h9c52;
sos_loop[0].somModel.sram_ptr[5][278]=3;
sos_loop[0].somModel.sram_dat[5][279][0]=96'h8583;
sos_loop[0].somModel.sram_ptr[5][279]=3;
sos_loop[0].somModel.sram_dat[5][280][0]=96'hf1e2;
sos_loop[0].somModel.sram_ptr[5][280]=3;
sos_loop[0].somModel.sram_dat[5][281][0]=96'hb68d;
sos_loop[0].somModel.sram_ptr[5][281]=3;
sos_loop[0].somModel.sram_dat[5][282][0]=96'h22c5;
sos_loop[0].somModel.sram_ptr[5][282]=3;
sos_loop[0].somModel.sram_dat[5][283][0]=96'h35a0;
sos_loop[0].somModel.sram_ptr[5][283]=3;
sos_loop[0].somModel.sram_dat[5][284][0]=96'hd202;
sos_loop[0].somModel.sram_ptr[5][284]=3;
sos_loop[0].somModel.sram_dat[5][285][0]=96'h87af;
sos_loop[0].somModel.sram_ptr[5][285]=3;
sos_loop[0].somModel.sram_dat[5][286][0]=96'hf3b0;
sos_loop[0].somModel.sram_ptr[5][286]=3;
sos_loop[0].somModel.sram_dat[5][287][0]=96'h646e;
sos_loop[0].somModel.sram_ptr[5][287]=3;
sos_loop[0].somModel.sram_dat[5][288][0]=96'h227e;
sos_loop[0].somModel.sram_ptr[5][288]=3;
sos_loop[0].somModel.sram_dat[5][289][0]=96'hdbb4;
sos_loop[0].somModel.sram_ptr[5][289]=3;
sos_loop[0].somModel.sram_dat[5][290][0]=96'h2830;
sos_loop[0].somModel.sram_ptr[5][290]=3;
sos_loop[0].somModel.sram_dat[5][291][0]=96'hf47;
sos_loop[0].somModel.sram_ptr[5][291]=3;
sos_loop[0].somModel.sram_dat[5][292][0]=96'h6e3a;
sos_loop[0].somModel.sram_ptr[5][292]=3;
sos_loop[0].somModel.sram_dat[5][293][0]=96'h13f3;
sos_loop[0].somModel.sram_ptr[5][293]=3;
sos_loop[0].somModel.sram_dat[5][294][0]=96'h4667;
sos_loop[0].somModel.sram_ptr[5][294]=3;
sos_loop[0].somModel.sram_dat[5][295][0]=96'h39b8;
sos_loop[0].somModel.sram_ptr[5][295]=3;
sos_loop[0].somModel.sram_dat[5][296][0]=96'h54e5;
sos_loop[0].somModel.sram_ptr[5][296]=3;
sos_loop[0].somModel.sram_dat[5][297][0]=96'h58ec;
sos_loop[0].somModel.sram_ptr[5][297]=3;
sos_loop[0].somModel.sram_dat[5][298][0]=96'h6869;
sos_loop[0].somModel.sram_ptr[5][298]=3;
sos_loop[0].somModel.sram_dat[5][299][0]=96'h6bbe;
sos_loop[0].somModel.sram_ptr[5][299]=3;
sos_loop[0].somModel.sram_dat[5][300][0]=96'h7815;
sos_loop[0].somModel.sram_ptr[5][300]=3;
sos_loop[0].somModel.sram_dat[5][301][0]=96'hd546;
sos_loop[0].somModel.sram_ptr[5][301]=3;
sos_loop[0].somModel.sram_dat[5][302][0]=96'h68ce;
sos_loop[0].somModel.sram_ptr[5][302]=3;
sos_loop[0].somModel.sram_dat[5][303][0]=96'hec8a;
sos_loop[0].somModel.sram_ptr[5][303]=3;
sos_loop[0].somModel.sram_dat[5][304][0]=96'hfb29;
sos_loop[0].somModel.sram_ptr[5][304]=3;
sos_loop[0].somModel.sram_dat[5][305][0]=96'hc7a;
sos_loop[0].somModel.sram_ptr[5][305]=3;
sos_loop[0].somModel.sram_dat[5][306][0]=96'h4760;
sos_loop[0].somModel.sram_ptr[5][306]=3;
sos_loop[0].somModel.sram_dat[5][307][0]=96'h34fc;
sos_loop[0].somModel.sram_ptr[5][307]=3;
sos_loop[0].somModel.sram_dat[5][308][0]=96'h7313;
sos_loop[0].somModel.sram_ptr[5][308]=3;
sos_loop[0].somModel.sram_dat[5][309][0]=96'ha699;
sos_loop[0].somModel.sram_ptr[5][309]=3;
sos_loop[0].somModel.sram_dat[5][310][0]=96'hd724;
sos_loop[0].somModel.sram_ptr[5][310]=3;
sos_loop[0].somModel.sram_dat[5][311][0]=96'hd427;
sos_loop[0].somModel.sram_ptr[5][311]=3;
sos_loop[0].somModel.sram_dat[5][312][0]=96'hefcd;
sos_loop[0].somModel.sram_ptr[5][312]=3;
sos_loop[0].somModel.sram_dat[5][313][0]=96'hf203;
sos_loop[0].somModel.sram_ptr[5][313]=3;
sos_loop[0].somModel.sram_dat[5][314][0]=96'h41da;
sos_loop[0].somModel.sram_ptr[5][314]=3;
sos_loop[0].somModel.sram_dat[5][315][0]=96'h390c;
sos_loop[0].somModel.sram_ptr[5][315]=3;
sos_loop[0].somModel.sram_dat[5][316][0]=96'h4b5a;
sos_loop[0].somModel.sram_ptr[5][316]=3;
sos_loop[0].somModel.sram_dat[5][317][0]=96'hc980;
sos_loop[0].somModel.sram_ptr[5][317]=3;
sos_loop[0].somModel.sram_dat[5][318][0]=96'hf62d;
sos_loop[0].somModel.sram_ptr[5][318]=3;
sos_loop[0].somModel.sram_dat[5][319][0]=96'h6fe6;
sos_loop[0].somModel.sram_ptr[5][319]=3;
sos_loop[0].somModel.sram_dat[5][320][0]=96'h8e36;
sos_loop[0].somModel.sram_ptr[5][320]=3;
sos_loop[0].somModel.sram_dat[5][321][0]=96'h32cc;
sos_loop[0].somModel.sram_ptr[5][321]=3;
sos_loop[0].somModel.sram_dat[5][322][0]=96'hab0e;
sos_loop[0].somModel.sram_ptr[5][322]=3;
sos_loop[0].somModel.sram_dat[5][323][0]=96'h87e8;
sos_loop[0].somModel.sram_ptr[5][323]=3;
sos_loop[0].somModel.sram_dat[5][324][0]=96'hc504;
sos_loop[0].somModel.sram_ptr[5][324]=3;
sos_loop[0].somModel.sram_dat[5][325][0]=96'h2a99;
sos_loop[0].somModel.sram_ptr[5][325]=3;
sos_loop[0].somModel.sram_dat[5][326][0]=96'h6e23;
sos_loop[0].somModel.sram_ptr[5][326]=3;
sos_loop[0].somModel.sram_dat[5][327][0]=96'h7936;
sos_loop[0].somModel.sram_ptr[5][327]=3;
sos_loop[0].somModel.sram_dat[5][328][0]=96'he3be;
sos_loop[0].somModel.sram_ptr[5][328]=3;
sos_loop[0].somModel.sram_dat[5][329][0]=96'h3d8c;
sos_loop[0].somModel.sram_ptr[5][329]=3;
sos_loop[0].somModel.sram_dat[5][330][0]=96'h689f;
sos_loop[0].somModel.sram_ptr[5][330]=3;
sos_loop[0].somModel.sram_dat[5][331][0]=96'hd3c9;
sos_loop[0].somModel.sram_ptr[5][331]=3;
sos_loop[0].somModel.sram_dat[5][332][0]=96'hcf80;
sos_loop[0].somModel.sram_ptr[5][332]=3;
sos_loop[0].somModel.sram_dat[5][333][0]=96'hc8b4;
sos_loop[0].somModel.sram_ptr[5][333]=3;
sos_loop[0].somModel.sram_dat[5][334][0]=96'h7438;
sos_loop[0].somModel.sram_ptr[5][334]=3;
sos_loop[0].somModel.sram_dat[5][335][0]=96'hd02d;
sos_loop[0].somModel.sram_ptr[5][335]=3;
sos_loop[0].somModel.sram_dat[5][336][0]=96'h5653;
sos_loop[0].somModel.sram_ptr[5][336]=3;
sos_loop[0].somModel.sram_dat[5][337][0]=96'h462a;
sos_loop[0].somModel.sram_ptr[5][337]=3;
sos_loop[0].somModel.sram_dat[5][338][0]=96'h79b6;
sos_loop[0].somModel.sram_ptr[5][338]=3;
sos_loop[0].somModel.sram_dat[5][339][0]=96'hff26;
sos_loop[0].somModel.sram_ptr[5][339]=3;
sos_loop[0].somModel.sram_dat[5][340][0]=96'hc9f8;
sos_loop[0].somModel.sram_ptr[5][340]=3;
sos_loop[0].somModel.sram_dat[5][341][0]=96'hc4de;
sos_loop[0].somModel.sram_ptr[5][341]=3;
sos_loop[0].somModel.sram_dat[5][342][0]=96'hfd4b;
sos_loop[0].somModel.sram_ptr[5][342]=3;
sos_loop[0].somModel.sram_dat[5][343][0]=96'h1cc0;
sos_loop[0].somModel.sram_ptr[5][343]=3;
sos_loop[0].somModel.sram_dat[5][344][0]=96'h3961;
sos_loop[0].somModel.sram_ptr[5][344]=3;
sos_loop[0].somModel.sram_dat[5][345][0]=96'hfac3;
sos_loop[0].somModel.sram_ptr[5][345]=3;
sos_loop[0].somModel.sram_dat[5][346][0]=96'h96b3;
sos_loop[0].somModel.sram_ptr[5][346]=3;
sos_loop[0].somModel.sram_dat[5][347][0]=96'h1d75;
sos_loop[0].somModel.sram_ptr[5][347]=3;
sos_loop[0].somModel.sram_dat[5][348][0]=96'hfeeb;
sos_loop[0].somModel.sram_ptr[5][348]=3;
sos_loop[0].somModel.sram_dat[5][349][0]=96'hd35;
sos_loop[0].somModel.sram_ptr[5][349]=3;
sos_loop[0].somModel.sram_dat[5][350][0]=96'hc987;
sos_loop[0].somModel.sram_ptr[5][350]=3;
sos_loop[0].somModel.sram_dat[5][351][0]=96'h3659;
sos_loop[0].somModel.sram_ptr[5][351]=3;
sos_loop[0].somModel.sram_dat[5][352][0]=96'hed9a;
sos_loop[0].somModel.sram_ptr[5][352]=3;
sos_loop[0].somModel.sram_dat[5][353][0]=96'ha77d;
sos_loop[0].somModel.sram_ptr[5][353]=3;
sos_loop[0].somModel.sram_dat[5][354][0]=96'hea;
sos_loop[0].somModel.sram_ptr[5][354]=3;
sos_loop[0].somModel.sram_dat[5][355][0]=96'h6d0c;
sos_loop[0].somModel.sram_ptr[5][355]=3;
sos_loop[0].somModel.sram_dat[5][356][0]=96'h5f79;
sos_loop[0].somModel.sram_ptr[5][356]=3;
sos_loop[0].somModel.sram_dat[5][357][0]=96'h3ab0;
sos_loop[0].somModel.sram_ptr[5][357]=3;
sos_loop[0].somModel.sram_dat[5][358][0]=96'h977e;
sos_loop[0].somModel.sram_ptr[5][358]=3;
sos_loop[0].somModel.sram_dat[5][359][0]=96'h3413;
sos_loop[0].somModel.sram_ptr[5][359]=3;
sos_loop[0].somModel.sram_dat[5][360][0]=96'h990c;
sos_loop[0].somModel.sram_ptr[5][360]=3;
sos_loop[0].somModel.sram_dat[5][361][0]=96'h530f;
sos_loop[0].somModel.sram_ptr[5][361]=3;
sos_loop[0].somModel.sram_dat[5][362][0]=96'h9949;
sos_loop[0].somModel.sram_ptr[5][362]=3;
sos_loop[0].somModel.sram_dat[5][363][0]=96'he132;
sos_loop[0].somModel.sram_ptr[5][363]=3;
sos_loop[0].somModel.sram_dat[5][364][0]=96'h47e1;
sos_loop[0].somModel.sram_ptr[5][364]=3;
sos_loop[0].somModel.sram_dat[5][365][0]=96'h77a2;
sos_loop[0].somModel.sram_ptr[5][365]=3;
sos_loop[0].somModel.sram_dat[5][366][0]=96'hb608;
sos_loop[0].somModel.sram_ptr[5][366]=3;
sos_loop[0].somModel.sram_dat[5][367][0]=96'ha7e7;
sos_loop[0].somModel.sram_ptr[5][367]=3;
sos_loop[0].somModel.sram_dat[5][368][0]=96'hd940;
sos_loop[0].somModel.sram_ptr[5][368]=3;
sos_loop[0].somModel.sram_dat[5][369][0]=96'hfb69;
sos_loop[0].somModel.sram_ptr[5][369]=3;
sos_loop[0].somModel.sram_dat[5][370][0]=96'h131c;
sos_loop[0].somModel.sram_ptr[5][370]=3;
sos_loop[0].somModel.sram_dat[5][371][0]=96'h5d26;
sos_loop[0].somModel.sram_ptr[5][371]=3;
sos_loop[0].somModel.sram_dat[5][372][0]=96'ha9cc;
sos_loop[0].somModel.sram_ptr[5][372]=3;
sos_loop[0].somModel.sram_dat[5][373][0]=96'h3677;
sos_loop[0].somModel.sram_ptr[5][373]=3;
sos_loop[0].somModel.sram_dat[5][374][0]=96'h4a66;
sos_loop[0].somModel.sram_ptr[5][374]=3;
sos_loop[0].somModel.sram_dat[5][375][0]=96'h9b09;
sos_loop[0].somModel.sram_ptr[5][375]=3;
sos_loop[0].somModel.sram_dat[5][376][0]=96'h3cea;
sos_loop[0].somModel.sram_ptr[5][376]=3;
sos_loop[0].somModel.sram_dat[5][377][0]=96'h4f86;
sos_loop[0].somModel.sram_ptr[5][377]=3;
sos_loop[0].somModel.sram_dat[5][378][0]=96'h5443;
sos_loop[0].somModel.sram_ptr[5][378]=3;
sos_loop[0].somModel.sram_dat[5][379][0]=96'hcc10;
sos_loop[0].somModel.sram_ptr[5][379]=3;
sos_loop[0].somModel.sram_dat[5][380][0]=96'ha83c;
sos_loop[0].somModel.sram_ptr[5][380]=3;
sos_loop[0].somModel.sram_dat[5][381][0]=96'h2399;
sos_loop[0].somModel.sram_ptr[5][381]=3;
sos_loop[0].somModel.sram_dat[5][382][0]=96'heed1;
sos_loop[0].somModel.sram_ptr[5][382]=3;
sos_loop[0].somModel.sram_dat[5][383][0]=96'h8b00;
sos_loop[0].somModel.sram_ptr[5][383]=3;
sos_loop[0].somModel.sram_dat[5][384][0]=96'hc875;
sos_loop[0].somModel.sram_ptr[5][384]=3;
sos_loop[0].somModel.sram_dat[5][385][0]=96'h30e5;
sos_loop[0].somModel.sram_ptr[5][385]=3;
sos_loop[0].somModel.sram_dat[5][386][0]=96'hc912;
sos_loop[0].somModel.sram_ptr[5][386]=3;
sos_loop[0].somModel.sram_dat[5][387][0]=96'h95c2;
sos_loop[0].somModel.sram_ptr[5][387]=3;
sos_loop[0].somModel.sram_dat[5][388][0]=96'hf263;
sos_loop[0].somModel.sram_ptr[5][388]=3;
sos_loop[0].somModel.sram_dat[5][389][0]=96'h5500;
sos_loop[0].somModel.sram_ptr[5][389]=3;
sos_loop[0].somModel.sram_dat[5][390][0]=96'h3863;
sos_loop[0].somModel.sram_ptr[5][390]=3;
sos_loop[0].somModel.sram_dat[5][391][0]=96'hda52;
sos_loop[0].somModel.sram_ptr[5][391]=3;
sos_loop[0].somModel.sram_dat[5][392][0]=96'h4a7f;
sos_loop[0].somModel.sram_ptr[5][392]=3;
sos_loop[0].somModel.sram_dat[5][393][0]=96'h31b;
sos_loop[0].somModel.sram_ptr[5][393]=3;
sos_loop[0].somModel.sram_dat[5][394][0]=96'h1bac;
sos_loop[0].somModel.sram_ptr[5][394]=3;
sos_loop[0].somModel.sram_dat[5][395][0]=96'h9b43;
sos_loop[0].somModel.sram_ptr[5][395]=3;
sos_loop[0].somModel.sram_dat[5][396][0]=96'ha30f;
sos_loop[0].somModel.sram_ptr[5][396]=3;
sos_loop[0].somModel.sram_dat[5][397][0]=96'hc88d;
sos_loop[0].somModel.sram_ptr[5][397]=3;
sos_loop[0].somModel.sram_dat[5][398][0]=96'h1146;
sos_loop[0].somModel.sram_ptr[5][398]=3;
sos_loop[0].somModel.sram_dat[5][399][0]=96'h33e3;
sos_loop[0].somModel.sram_ptr[5][399]=3;
sos_loop[0].somModel.sram_dat[5][400][0]=96'hd222;
sos_loop[0].somModel.sram_ptr[5][400]=3;
sos_loop[0].somModel.sram_dat[5][401][0]=96'hbf0a;
sos_loop[0].somModel.sram_ptr[5][401]=3;
sos_loop[0].somModel.sram_dat[5][402][0]=96'h8d89;
sos_loop[0].somModel.sram_ptr[5][402]=3;
sos_loop[0].somModel.sram_dat[5][403][0]=96'h24f0;
sos_loop[0].somModel.sram_ptr[5][403]=3;
sos_loop[0].somModel.sram_dat[5][404][0]=96'he2e;
sos_loop[0].somModel.sram_ptr[5][404]=3;
sos_loop[0].somModel.sram_dat[5][405][0]=96'hd40c;
sos_loop[0].somModel.sram_ptr[5][405]=3;
sos_loop[0].somModel.sram_dat[5][406][0]=96'h2570;
sos_loop[0].somModel.sram_ptr[5][406]=3;
sos_loop[0].somModel.sram_dat[5][407][0]=96'h2acc;
sos_loop[0].somModel.sram_ptr[5][407]=3;
sos_loop[0].somModel.sram_dat[5][408][0]=96'h3dc1;
sos_loop[0].somModel.sram_ptr[5][408]=3;
sos_loop[0].somModel.sram_dat[5][409][0]=96'h5b5b;
sos_loop[0].somModel.sram_ptr[5][409]=3;
sos_loop[0].somModel.sram_dat[5][410][0]=96'h4198;
sos_loop[0].somModel.sram_ptr[5][410]=3;
sos_loop[0].somModel.sram_dat[5][411][0]=96'h8e6d;
sos_loop[0].somModel.sram_ptr[5][411]=3;
sos_loop[0].somModel.sram_dat[5][412][0]=96'h12a8;
sos_loop[0].somModel.sram_ptr[5][412]=3;
sos_loop[0].somModel.sram_dat[5][413][0]=96'hfd89;
sos_loop[0].somModel.sram_ptr[5][413]=3;
sos_loop[0].somModel.sram_dat[5][414][0]=96'h2577;
sos_loop[0].somModel.sram_ptr[5][414]=3;
sos_loop[0].somModel.sram_dat[5][415][0]=96'h3edf;
sos_loop[0].somModel.sram_ptr[5][415]=3;
sos_loop[0].somModel.sram_dat[5][416][0]=96'h6331;
sos_loop[0].somModel.sram_ptr[5][416]=3;
sos_loop[0].somModel.sram_dat[5][417][0]=96'h4747;
sos_loop[0].somModel.sram_ptr[5][417]=3;
sos_loop[0].somModel.sram_dat[5][418][0]=96'h2327;
sos_loop[0].somModel.sram_ptr[5][418]=3;
sos_loop[0].somModel.sram_dat[5][419][0]=96'h4c09;
sos_loop[0].somModel.sram_ptr[5][419]=3;
sos_loop[0].somModel.sram_dat[5][420][0]=96'h1a17;
sos_loop[0].somModel.sram_ptr[5][420]=3;
sos_loop[0].somModel.sram_dat[5][421][0]=96'ha395;
sos_loop[0].somModel.sram_ptr[5][421]=3;
sos_loop[0].somModel.sram_dat[5][422][0]=96'hc94;
sos_loop[0].somModel.sram_ptr[5][422]=3;
sos_loop[0].somModel.sram_dat[5][423][0]=96'h174;
sos_loop[0].somModel.sram_ptr[5][423]=3;
sos_loop[0].somModel.sram_dat[5][424][0]=96'h212e;
sos_loop[0].somModel.sram_ptr[5][424]=3;
sos_loop[0].somModel.sram_dat[5][425][0]=96'h80ab;
sos_loop[0].somModel.sram_ptr[5][425]=3;
sos_loop[0].somModel.sram_dat[5][426][0]=96'ha361;
sos_loop[0].somModel.sram_ptr[5][426]=3;
sos_loop[0].somModel.sram_dat[5][427][0]=96'hfbf6;
sos_loop[0].somModel.sram_ptr[5][427]=3;
sos_loop[0].somModel.sram_dat[5][428][0]=96'hd291;
sos_loop[0].somModel.sram_ptr[5][428]=3;
sos_loop[0].somModel.sram_dat[5][429][0]=96'h81bf;
sos_loop[0].somModel.sram_ptr[5][429]=3;
sos_loop[0].somModel.sram_dat[5][430][0]=96'hc9e;
sos_loop[0].somModel.sram_ptr[5][430]=3;
sos_loop[0].somModel.sram_dat[5][431][0]=96'he846;
sos_loop[0].somModel.sram_ptr[5][431]=3;
sos_loop[0].somModel.sram_dat[5][432][0]=96'hd5c;
sos_loop[0].somModel.sram_ptr[5][432]=3;
sos_loop[0].somModel.sram_dat[5][433][0]=96'hce2a;
sos_loop[0].somModel.sram_ptr[5][433]=3;
sos_loop[0].somModel.sram_dat[5][434][0]=96'hfa53;
sos_loop[0].somModel.sram_ptr[5][434]=3;
sos_loop[0].somModel.sram_dat[5][435][0]=96'h4afe;
sos_loop[0].somModel.sram_ptr[5][435]=3;
sos_loop[0].somModel.sram_dat[5][436][0]=96'h215d;
sos_loop[0].somModel.sram_ptr[5][436]=3;
sos_loop[0].somModel.sram_dat[5][437][0]=96'ha8f9;
sos_loop[0].somModel.sram_ptr[5][437]=3;
sos_loop[0].somModel.sram_dat[5][438][0]=96'h9fff;
sos_loop[0].somModel.sram_ptr[5][438]=3;
sos_loop[0].somModel.sram_dat[5][439][0]=96'h539d;
sos_loop[0].somModel.sram_ptr[5][439]=3;
sos_loop[0].somModel.sram_dat[5][440][0]=96'h2c1e;
sos_loop[0].somModel.sram_ptr[5][440]=3;
sos_loop[0].somModel.sram_dat[5][441][0]=96'h3ea8;
sos_loop[0].somModel.sram_ptr[5][441]=3;
sos_loop[0].somModel.sram_dat[5][442][0]=96'h8d4c;
sos_loop[0].somModel.sram_ptr[5][442]=3;
sos_loop[0].somModel.sram_dat[5][443][0]=96'h9c5c;
sos_loop[0].somModel.sram_ptr[5][443]=3;
sos_loop[0].somModel.sram_dat[5][444][0]=96'hdb37;
sos_loop[0].somModel.sram_ptr[5][444]=3;
sos_loop[0].somModel.sram_dat[5][445][0]=96'ha769;
sos_loop[0].somModel.sram_ptr[5][445]=3;
sos_loop[0].somModel.sram_dat[5][446][0]=96'h1c12;
sos_loop[0].somModel.sram_ptr[5][446]=3;
sos_loop[0].somModel.sram_dat[5][447][0]=96'h42e3;
sos_loop[0].somModel.sram_ptr[5][447]=3;
sos_loop[0].somModel.sram_dat[5][448][0]=96'hc8ca;
sos_loop[0].somModel.sram_ptr[5][448]=3;
sos_loop[0].somModel.sram_dat[5][449][0]=96'hacf8;
sos_loop[0].somModel.sram_ptr[5][449]=3;
sos_loop[0].somModel.sram_dat[5][450][0]=96'hf770;
sos_loop[0].somModel.sram_ptr[5][450]=3;
sos_loop[0].somModel.sram_dat[5][451][0]=96'h57ff;
sos_loop[0].somModel.sram_ptr[5][451]=3;
sos_loop[0].somModel.sram_dat[5][452][0]=96'h6a40;
sos_loop[0].somModel.sram_ptr[5][452]=3;
sos_loop[0].somModel.sram_dat[5][453][0]=96'h6579;
sos_loop[0].somModel.sram_ptr[5][453]=3;
sos_loop[0].somModel.sram_dat[5][454][0]=96'h499e;
sos_loop[0].somModel.sram_ptr[5][454]=3;
sos_loop[0].somModel.sram_dat[5][455][0]=96'h27a1;
sos_loop[0].somModel.sram_ptr[5][455]=3;
sos_loop[0].somModel.sram_dat[5][456][0]=96'h9123;
sos_loop[0].somModel.sram_ptr[5][456]=3;
sos_loop[0].somModel.sram_dat[5][457][0]=96'ha641;
sos_loop[0].somModel.sram_ptr[5][457]=3;
sos_loop[0].somModel.sram_dat[5][458][0]=96'h80db;
sos_loop[0].somModel.sram_ptr[5][458]=3;
sos_loop[0].somModel.sram_dat[5][459][0]=96'hcbf3;
sos_loop[0].somModel.sram_ptr[5][459]=3;
sos_loop[0].somModel.sram_dat[5][460][0]=96'ha9a5;
sos_loop[0].somModel.sram_ptr[5][460]=3;
sos_loop[0].somModel.sram_dat[5][461][0]=96'h3824;
sos_loop[0].somModel.sram_ptr[5][461]=3;
sos_loop[0].somModel.sram_dat[5][462][0]=96'hc25d;
sos_loop[0].somModel.sram_ptr[5][462]=3;
sos_loop[0].somModel.sram_dat[5][463][0]=96'hd240;
sos_loop[0].somModel.sram_ptr[5][463]=3;
sos_loop[0].somModel.sram_dat[5][464][0]=96'hbebd;
sos_loop[0].somModel.sram_ptr[5][464]=3;
sos_loop[0].somModel.sram_dat[5][465][0]=96'he5fc;
sos_loop[0].somModel.sram_ptr[5][465]=3;
sos_loop[0].somModel.sram_dat[5][466][0]=96'h7e08;
sos_loop[0].somModel.sram_ptr[5][466]=3;
sos_loop[0].somModel.sram_dat[5][467][0]=96'h6999;
sos_loop[0].somModel.sram_ptr[5][467]=3;
sos_loop[0].somModel.sram_dat[5][468][0]=96'ha30b;
sos_loop[0].somModel.sram_ptr[5][468]=3;
sos_loop[0].somModel.sram_dat[5][469][0]=96'hb086;
sos_loop[0].somModel.sram_ptr[5][469]=3;
sos_loop[0].somModel.sram_dat[5][470][0]=96'h2c3e;
sos_loop[0].somModel.sram_ptr[5][470]=3;
sos_loop[0].somModel.sram_dat[5][471][0]=96'he232;
sos_loop[0].somModel.sram_ptr[5][471]=3;
sos_loop[0].somModel.sram_dat[5][472][0]=96'hc378;
sos_loop[0].somModel.sram_ptr[5][472]=3;
sos_loop[0].somModel.sram_dat[5][473][0]=96'hb14c;
sos_loop[0].somModel.sram_ptr[5][473]=3;
sos_loop[0].somModel.sram_dat[5][474][0]=96'h2bb7;
sos_loop[0].somModel.sram_ptr[5][474]=3;
sos_loop[0].somModel.sram_dat[5][475][0]=96'hd28;
sos_loop[0].somModel.sram_ptr[5][475]=3;
sos_loop[0].somModel.sram_dat[5][476][0]=96'hb678;
sos_loop[0].somModel.sram_ptr[5][476]=3;
sos_loop[0].somModel.sram_dat[5][477][0]=96'ha845;
sos_loop[0].somModel.sram_ptr[5][477]=3;
sos_loop[0].somModel.sram_dat[5][478][0]=96'hc805;
sos_loop[0].somModel.sram_ptr[5][478]=3;
sos_loop[0].somModel.sram_dat[5][479][0]=96'hf905;
sos_loop[0].somModel.sram_ptr[5][479]=3;
sos_loop[0].somModel.sram_dat[5][480][0]=96'h5909;
sos_loop[0].somModel.sram_ptr[5][480]=3;
sos_loop[0].somModel.sram_dat[5][481][0]=96'h1850;
sos_loop[0].somModel.sram_ptr[5][481]=3;
sos_loop[0].somModel.sram_dat[5][482][0]=96'h3708;
sos_loop[0].somModel.sram_ptr[5][482]=3;
sos_loop[0].somModel.sram_dat[5][483][0]=96'h3bb1;
sos_loop[0].somModel.sram_ptr[5][483]=3;
sos_loop[0].somModel.sram_dat[5][484][0]=96'hfe35;
sos_loop[0].somModel.sram_ptr[5][484]=3;
sos_loop[0].somModel.sram_dat[5][485][0]=96'h3010;
sos_loop[0].somModel.sram_ptr[5][485]=3;
sos_loop[0].somModel.sram_dat[5][486][0]=96'h222f;
sos_loop[0].somModel.sram_ptr[5][486]=3;
sos_loop[0].somModel.sram_dat[5][487][0]=96'h56fa;
sos_loop[0].somModel.sram_ptr[5][487]=3;
sos_loop[0].somModel.sram_dat[5][488][0]=96'h3023;
sos_loop[0].somModel.sram_ptr[5][488]=3;
sos_loop[0].somModel.sram_dat[5][489][0]=96'hde51;
sos_loop[0].somModel.sram_ptr[5][489]=3;
sos_loop[0].somModel.sram_dat[5][490][0]=96'h9900;
sos_loop[0].somModel.sram_ptr[5][490]=3;
sos_loop[0].somModel.sram_dat[5][491][0]=96'h7b27;
sos_loop[0].somModel.sram_ptr[5][491]=3;
sos_loop[0].somModel.sram_dat[5][492][0]=96'ha678;
sos_loop[0].somModel.sram_ptr[5][492]=3;
sos_loop[0].somModel.sram_dat[5][493][0]=96'h4ff3;
sos_loop[0].somModel.sram_ptr[5][493]=3;
sos_loop[0].somModel.sram_dat[5][494][0]=96'h95fc;
sos_loop[0].somModel.sram_ptr[5][494]=3;
sos_loop[0].somModel.sram_dat[5][495][0]=96'h8d2c;
sos_loop[0].somModel.sram_ptr[5][495]=3;
sos_loop[0].somModel.sram_dat[5][496][0]=96'h8a9e;
sos_loop[0].somModel.sram_ptr[5][496]=3;
sos_loop[0].somModel.sram_dat[5][497][0]=96'heef;
sos_loop[0].somModel.sram_ptr[5][497]=3;
sos_loop[0].somModel.sram_dat[5][498][0]=96'hd8e7;
sos_loop[0].somModel.sram_ptr[5][498]=3;
sos_loop[0].somModel.sram_dat[5][499][0]=96'ha7e;
sos_loop[0].somModel.sram_ptr[5][499]=3;
sos_loop[0].somModel.sram_dat[5][500][0]=96'h19a1;
sos_loop[0].somModel.sram_ptr[5][500]=3;
sos_loop[0].somModel.sram_dat[5][501][0]=96'hec33;
sos_loop[0].somModel.sram_ptr[5][501]=3;
sos_loop[0].somModel.sram_dat[5][502][0]=96'ha05a;
sos_loop[0].somModel.sram_ptr[5][502]=3;
sos_loop[0].somModel.sram_dat[5][503][0]=96'h7046;
sos_loop[0].somModel.sram_ptr[5][503]=3;
sos_loop[0].somModel.sram_dat[5][504][0]=96'h2ea1;
sos_loop[0].somModel.sram_ptr[5][504]=3;
sos_loop[0].somModel.sram_dat[5][505][0]=96'h9bf1;
sos_loop[0].somModel.sram_ptr[5][505]=3;
sos_loop[0].somModel.sram_dat[5][506][0]=96'hac89;
sos_loop[0].somModel.sram_ptr[5][506]=3;
sos_loop[0].somModel.sram_dat[5][507][0]=96'h1572;
sos_loop[0].somModel.sram_ptr[5][507]=3;
sos_loop[0].somModel.sram_dat[5][508][0]=96'h1b4c;
sos_loop[0].somModel.sram_ptr[5][508]=3;
sos_loop[0].somModel.sram_dat[5][509][0]=96'h66b0;
sos_loop[0].somModel.sram_ptr[5][509]=3;
sos_loop[0].somModel.sram_dat[5][510][0]=96'h46e;
sos_loop[0].somModel.sram_ptr[5][510]=3;
sos_loop[0].somModel.sram_dat[5][511][0]=96'hf521;
sos_loop[0].somModel.sram_ptr[5][511]=3;
sos_loop[0].somModel.sram_dat[5][512][0]=96'h7fed;
sos_loop[0].somModel.sram_ptr[5][512]=3;
sos_loop[0].somModel.sram_dat[5][513][0]=96'ha538;
sos_loop[0].somModel.sram_ptr[5][513]=3;
sos_loop[0].somModel.sram_dat[5][514][0]=96'h721d;
sos_loop[0].somModel.sram_ptr[5][514]=3;
sos_loop[0].somModel.sram_dat[5][515][0]=96'h1f85;
sos_loop[0].somModel.sram_ptr[5][515]=3;
sos_loop[0].somModel.sram_dat[5][516][0]=96'hddcf;
sos_loop[0].somModel.sram_ptr[5][516]=3;
sos_loop[0].somModel.sram_dat[5][517][0]=96'h923c;
sos_loop[0].somModel.sram_ptr[5][517]=3;
sos_loop[0].somModel.sram_dat[5][518][0]=96'h5be3;
sos_loop[0].somModel.sram_ptr[5][518]=3;
sos_loop[0].somModel.sram_dat[5][519][0]=96'hc41c;
sos_loop[0].somModel.sram_ptr[5][519]=3;
sos_loop[0].somModel.sram_dat[5][520][0]=96'he73;
sos_loop[0].somModel.sram_ptr[5][520]=3;
sos_loop[0].somModel.sram_dat[5][521][0]=96'h4046;
sos_loop[0].somModel.sram_ptr[5][521]=3;
sos_loop[0].somModel.sram_dat[5][522][0]=96'h8109;
sos_loop[0].somModel.sram_ptr[5][522]=3;
sos_loop[0].somModel.sram_dat[5][523][0]=96'h966e;
sos_loop[0].somModel.sram_ptr[5][523]=3;
sos_loop[0].somModel.sram_dat[5][524][0]=96'he61a;
sos_loop[0].somModel.sram_ptr[5][524]=3;
sos_loop[0].somModel.sram_dat[5][525][0]=96'h7975;
sos_loop[0].somModel.sram_ptr[5][525]=3;
sos_loop[0].somModel.sram_dat[5][526][0]=96'hd88c;
sos_loop[0].somModel.sram_ptr[5][526]=3;
sos_loop[0].somModel.sram_dat[5][527][0]=96'h645a;
sos_loop[0].somModel.sram_ptr[5][527]=3;
sos_loop[0].somModel.sram_dat[5][528][0]=96'h87d2;
sos_loop[0].somModel.sram_ptr[5][528]=3;
sos_loop[0].somModel.sram_dat[5][529][0]=96'h619d;
sos_loop[0].somModel.sram_ptr[5][529]=3;
sos_loop[0].somModel.sram_dat[5][530][0]=96'h93fc;
sos_loop[0].somModel.sram_ptr[5][530]=3;
sos_loop[0].somModel.sram_dat[5][531][0]=96'h1d1b;
sos_loop[0].somModel.sram_ptr[5][531]=3;
sos_loop[0].somModel.sram_dat[5][532][0]=96'he191;
sos_loop[0].somModel.sram_ptr[5][532]=3;
sos_loop[0].somModel.sram_dat[5][533][0]=96'h8160;
sos_loop[0].somModel.sram_ptr[5][533]=3;
sos_loop[0].somModel.sram_dat[5][534][0]=96'hfd5e;
sos_loop[0].somModel.sram_ptr[5][534]=3;
sos_loop[0].somModel.sram_dat[5][535][0]=96'had9e;
sos_loop[0].somModel.sram_ptr[5][535]=3;
sos_loop[0].somModel.sram_dat[5][536][0]=96'he6bc;
sos_loop[0].somModel.sram_ptr[5][536]=3;
sos_loop[0].somModel.sram_dat[5][537][0]=96'h9199;
sos_loop[0].somModel.sram_ptr[5][537]=3;
sos_loop[0].somModel.sram_dat[5][538][0]=96'hffde;
sos_loop[0].somModel.sram_ptr[5][538]=3;
sos_loop[0].somModel.sram_dat[5][539][0]=96'h6c77;
sos_loop[0].somModel.sram_ptr[5][539]=3;
sos_loop[0].somModel.sram_dat[5][540][0]=96'h4d6c;
sos_loop[0].somModel.sram_ptr[5][540]=3;
sos_loop[0].somModel.sram_dat[5][541][0]=96'hd10a;
sos_loop[0].somModel.sram_ptr[5][541]=3;
sos_loop[0].somModel.sram_dat[5][542][0]=96'he977;
sos_loop[0].somModel.sram_ptr[5][542]=3;
sos_loop[0].somModel.sram_dat[5][543][0]=96'h4135;
sos_loop[0].somModel.sram_ptr[5][543]=3;
sos_loop[0].somModel.sram_dat[5][544][0]=96'hbcb9;
sos_loop[0].somModel.sram_ptr[5][544]=3;
sos_loop[0].somModel.sram_dat[5][545][0]=96'ha3ed;
sos_loop[0].somModel.sram_ptr[5][545]=3;
sos_loop[0].somModel.sram_dat[5][546][0]=96'h81ec;
sos_loop[0].somModel.sram_ptr[5][546]=3;
sos_loop[0].somModel.sram_dat[5][547][0]=96'h40f1;
sos_loop[0].somModel.sram_ptr[5][547]=3;
sos_loop[0].somModel.sram_dat[5][548][0]=96'he12e;
sos_loop[0].somModel.sram_ptr[5][548]=3;
sos_loop[0].somModel.sram_dat[5][549][0]=96'h8bd3;
sos_loop[0].somModel.sram_ptr[5][549]=3;
sos_loop[0].somModel.sram_dat[5][550][0]=96'h5de;
sos_loop[0].somModel.sram_ptr[5][550]=3;
sos_loop[0].somModel.sram_dat[5][551][0]=96'h852e;
sos_loop[0].somModel.sram_ptr[5][551]=3;
sos_loop[0].somModel.sram_dat[5][552][0]=96'h89be;
sos_loop[0].somModel.sram_ptr[5][552]=3;
sos_loop[0].somModel.sram_dat[5][553][0]=96'h9c0c;
sos_loop[0].somModel.sram_ptr[5][553]=3;
sos_loop[0].somModel.sram_dat[5][554][0]=96'h58fb;
sos_loop[0].somModel.sram_ptr[5][554]=3;
sos_loop[0].somModel.sram_dat[5][555][0]=96'haa88;
sos_loop[0].somModel.sram_ptr[5][555]=3;
sos_loop[0].somModel.sram_dat[5][556][0]=96'hb6f4;
sos_loop[0].somModel.sram_ptr[5][556]=3;
sos_loop[0].somModel.sram_dat[5][557][0]=96'h5206;
sos_loop[0].somModel.sram_ptr[5][557]=3;
sos_loop[0].somModel.sram_dat[5][558][0]=96'h6efd;
sos_loop[0].somModel.sram_ptr[5][558]=3;
sos_loop[0].somModel.sram_dat[5][559][0]=96'h432b;
sos_loop[0].somModel.sram_ptr[5][559]=3;
sos_loop[0].somModel.sram_dat[5][560][0]=96'h715e;
sos_loop[0].somModel.sram_ptr[5][560]=3;
sos_loop[0].somModel.sram_dat[5][561][0]=96'h633;
sos_loop[0].somModel.sram_ptr[5][561]=3;
sos_loop[0].somModel.sram_dat[5][562][0]=96'h9f03;
sos_loop[0].somModel.sram_ptr[5][562]=3;
sos_loop[0].somModel.sram_dat[5][563][0]=96'hed63;
sos_loop[0].somModel.sram_ptr[5][563]=3;
sos_loop[0].somModel.sram_dat[5][564][0]=96'h7a86;
sos_loop[0].somModel.sram_ptr[5][564]=3;
sos_loop[0].somModel.sram_dat[5][565][0]=96'h8df8;
sos_loop[0].somModel.sram_ptr[5][565]=3;
sos_loop[0].somModel.sram_dat[5][566][0]=96'h4007;
sos_loop[0].somModel.sram_ptr[5][566]=3;
sos_loop[0].somModel.sram_dat[5][567][0]=96'hdb34;
sos_loop[0].somModel.sram_ptr[5][567]=3;
sos_loop[0].somModel.sram_dat[5][568][0]=96'h7aa9;
sos_loop[0].somModel.sram_ptr[5][568]=3;
sos_loop[0].somModel.sram_dat[5][569][0]=96'h74d0;
sos_loop[0].somModel.sram_ptr[5][569]=3;
sos_loop[0].somModel.sram_dat[5][570][0]=96'hc8a5;
sos_loop[0].somModel.sram_ptr[5][570]=3;
sos_loop[0].somModel.sram_dat[5][571][0]=96'h2c9d;
sos_loop[0].somModel.sram_ptr[5][571]=3;
sos_loop[0].somModel.sram_dat[5][572][0]=96'h7b79;
sos_loop[0].somModel.sram_ptr[5][572]=3;
sos_loop[0].somModel.sram_dat[5][573][0]=96'hf1d6;
sos_loop[0].somModel.sram_ptr[5][573]=3;
sos_loop[0].somModel.sram_dat[5][574][0]=96'h8452;
sos_loop[0].somModel.sram_ptr[5][574]=3;
sos_loop[0].somModel.sram_dat[5][575][0]=96'ha758;
sos_loop[0].somModel.sram_ptr[5][575]=3;
sos_loop[0].somModel.sram_dat[5][576][0]=96'hc377;
sos_loop[0].somModel.sram_ptr[5][576]=3;
sos_loop[0].somModel.sram_dat[5][577][0]=96'h9a0a;
sos_loop[0].somModel.sram_ptr[5][577]=3;
sos_loop[0].somModel.sram_dat[5][578][0]=96'h51a0;
sos_loop[0].somModel.sram_ptr[5][578]=3;
sos_loop[0].somModel.sram_dat[5][579][0]=96'he2f5;
sos_loop[0].somModel.sram_ptr[5][579]=3;
sos_loop[0].somModel.sram_dat[5][580][0]=96'hebd0;
sos_loop[0].somModel.sram_ptr[5][580]=3;
sos_loop[0].somModel.sram_dat[5][581][0]=96'hbba;
sos_loop[0].somModel.sram_ptr[5][581]=3;
sos_loop[0].somModel.sram_dat[5][582][0]=96'h495a;
sos_loop[0].somModel.sram_ptr[5][582]=3;
sos_loop[0].somModel.sram_dat[5][583][0]=96'h84ac;
sos_loop[0].somModel.sram_ptr[5][583]=3;
sos_loop[0].somModel.sram_dat[5][584][0]=96'hd77;
sos_loop[0].somModel.sram_ptr[5][584]=3;
sos_loop[0].somModel.sram_dat[5][585][0]=96'hceef;
sos_loop[0].somModel.sram_ptr[5][585]=3;
sos_loop[0].somModel.sram_dat[5][586][0]=96'hbb05;
sos_loop[0].somModel.sram_ptr[5][586]=3;
sos_loop[0].somModel.sram_dat[5][587][0]=96'h7e66;
sos_loop[0].somModel.sram_ptr[5][587]=3;
sos_loop[0].somModel.sram_dat[5][588][0]=96'h6e53;
sos_loop[0].somModel.sram_ptr[5][588]=3;
sos_loop[0].somModel.sram_dat[5][589][0]=96'h9083;
sos_loop[0].somModel.sram_ptr[5][589]=3;
sos_loop[0].somModel.sram_dat[5][590][0]=96'h48cc;
sos_loop[0].somModel.sram_ptr[5][590]=3;
sos_loop[0].somModel.sram_dat[5][591][0]=96'h8be5;
sos_loop[0].somModel.sram_ptr[5][591]=3;
sos_loop[0].somModel.sram_dat[5][592][0]=96'h5f88;
sos_loop[0].somModel.sram_ptr[5][592]=3;
sos_loop[0].somModel.sram_dat[5][593][0]=96'h68a8;
sos_loop[0].somModel.sram_ptr[5][593]=3;
sos_loop[0].somModel.sram_dat[5][594][0]=96'hc805;
sos_loop[0].somModel.sram_ptr[5][594]=3;
sos_loop[0].somModel.sram_dat[5][595][0]=96'h9ecf;
sos_loop[0].somModel.sram_ptr[5][595]=3;
sos_loop[0].somModel.sram_dat[5][596][0]=96'hd5f0;
sos_loop[0].somModel.sram_ptr[5][596]=3;
sos_loop[0].somModel.sram_dat[5][597][0]=96'h1cfc;
sos_loop[0].somModel.sram_ptr[5][597]=3;
sos_loop[0].somModel.sram_dat[5][598][0]=96'hc265;
sos_loop[0].somModel.sram_ptr[5][598]=3;
sos_loop[0].somModel.sram_dat[5][599][0]=96'hd9b4;
sos_loop[0].somModel.sram_ptr[5][599]=3;
sos_loop[0].somModel.sram_dat[5][600][0]=96'h5053;
sos_loop[0].somModel.sram_ptr[5][600]=3;
sos_loop[0].somModel.sram_dat[5][601][0]=96'h6860;
sos_loop[0].somModel.sram_ptr[5][601]=3;
sos_loop[0].somModel.sram_dat[5][602][0]=96'h39a;
sos_loop[0].somModel.sram_ptr[5][602]=3;
sos_loop[0].somModel.sram_dat[5][603][0]=96'hbb6c;
sos_loop[0].somModel.sram_ptr[5][603]=3;
sos_loop[0].somModel.sram_dat[5][604][0]=96'h210c;
sos_loop[0].somModel.sram_ptr[5][604]=3;
sos_loop[0].somModel.sram_dat[5][605][0]=96'h6980;
sos_loop[0].somModel.sram_ptr[5][605]=3;
sos_loop[0].somModel.sram_dat[5][606][0]=96'ha25d;
sos_loop[0].somModel.sram_ptr[5][606]=3;
sos_loop[0].somModel.sram_dat[5][607][0]=96'h9aec;
sos_loop[0].somModel.sram_ptr[5][607]=3;
sos_loop[0].somModel.sram_dat[5][608][0]=96'hb8c5;
sos_loop[0].somModel.sram_ptr[5][608]=3;
sos_loop[0].somModel.sram_dat[5][609][0]=96'ha45b;
sos_loop[0].somModel.sram_ptr[5][609]=3;
sos_loop[0].somModel.sram_dat[5][610][0]=96'h1bfb;
sos_loop[0].somModel.sram_ptr[5][610]=3;
sos_loop[0].somModel.sram_dat[5][611][0]=96'h58d3;
sos_loop[0].somModel.sram_ptr[5][611]=3;
sos_loop[0].somModel.sram_dat[5][612][0]=96'he69;
sos_loop[0].somModel.sram_ptr[5][612]=3;
sos_loop[0].somModel.sram_dat[5][613][0]=96'h2820;
sos_loop[0].somModel.sram_ptr[5][613]=3;
sos_loop[0].somModel.sram_dat[5][614][0]=96'h4054;
sos_loop[0].somModel.sram_ptr[5][614]=3;
sos_loop[0].somModel.sram_dat[5][615][0]=96'hb2e2;
sos_loop[0].somModel.sram_ptr[5][615]=3;
sos_loop[0].somModel.sram_dat[5][616][0]=96'h316;
sos_loop[0].somModel.sram_ptr[5][616]=3;
sos_loop[0].somModel.sram_dat[5][617][0]=96'h7aa9;
sos_loop[0].somModel.sram_ptr[5][617]=3;
sos_loop[0].somModel.sram_dat[5][618][0]=96'h10a8;
sos_loop[0].somModel.sram_ptr[5][618]=3;
sos_loop[0].somModel.sram_dat[5][619][0]=96'he18a;
sos_loop[0].somModel.sram_ptr[5][619]=3;
sos_loop[0].somModel.sram_dat[5][620][0]=96'hab13;
sos_loop[0].somModel.sram_ptr[5][620]=3;
sos_loop[0].somModel.sram_dat[5][621][0]=96'hf1d1;
sos_loop[0].somModel.sram_ptr[5][621]=3;
sos_loop[0].somModel.sram_dat[5][622][0]=96'h14f2;
sos_loop[0].somModel.sram_ptr[5][622]=3;
sos_loop[0].somModel.sram_dat[5][623][0]=96'h6822;
sos_loop[0].somModel.sram_ptr[5][623]=3;
sos_loop[0].somModel.sram_dat[5][624][0]=96'h4228;
sos_loop[0].somModel.sram_ptr[5][624]=3;
sos_loop[0].somModel.sram_dat[5][625][0]=96'h81e5;
sos_loop[0].somModel.sram_ptr[5][625]=3;
sos_loop[0].somModel.sram_dat[5][626][0]=96'h6203;
sos_loop[0].somModel.sram_ptr[5][626]=3;
sos_loop[0].somModel.sram_dat[5][627][0]=96'h48b2;
sos_loop[0].somModel.sram_ptr[5][627]=3;
sos_loop[0].somModel.sram_dat[5][628][0]=96'h7b40;
sos_loop[0].somModel.sram_ptr[5][628]=3;
sos_loop[0].somModel.sram_dat[5][629][0]=96'hf692;
sos_loop[0].somModel.sram_ptr[5][629]=3;
sos_loop[0].somModel.sram_dat[5][630][0]=96'hab7e;
sos_loop[0].somModel.sram_ptr[5][630]=3;
sos_loop[0].somModel.sram_dat[5][631][0]=96'hce0c;
sos_loop[0].somModel.sram_ptr[5][631]=3;
sos_loop[0].somModel.sram_dat[5][632][0]=96'ha40b;
sos_loop[0].somModel.sram_ptr[5][632]=3;
sos_loop[0].somModel.sram_dat[5][633][0]=96'h4636;
sos_loop[0].somModel.sram_ptr[5][633]=3;
sos_loop[0].somModel.sram_dat[5][634][0]=96'h3aee;
sos_loop[0].somModel.sram_ptr[5][634]=3;
sos_loop[0].somModel.sram_dat[5][635][0]=96'hef6c;
sos_loop[0].somModel.sram_ptr[5][635]=3;
sos_loop[0].somModel.sram_dat[5][636][0]=96'h928f;
sos_loop[0].somModel.sram_ptr[5][636]=3;
sos_loop[0].somModel.sram_dat[5][637][0]=96'hd60f;
sos_loop[0].somModel.sram_ptr[5][637]=3;
sos_loop[0].somModel.sram_dat[5][638][0]=96'hbd68;
sos_loop[0].somModel.sram_ptr[5][638]=3;
sos_loop[0].somModel.sram_dat[5][639][0]=96'h30c9;
sos_loop[0].somModel.sram_ptr[5][639]=3;
sos_loop[0].somModel.sram_dat[5][640][0]=96'hcbd2;
sos_loop[0].somModel.sram_ptr[5][640]=3;
sos_loop[0].somModel.sram_dat[5][641][0]=96'hd53c;
sos_loop[0].somModel.sram_ptr[5][641]=3;
sos_loop[0].somModel.sram_dat[5][642][0]=96'h1685;
sos_loop[0].somModel.sram_ptr[5][642]=3;
sos_loop[0].somModel.sram_dat[5][643][0]=96'h2195;
sos_loop[0].somModel.sram_ptr[5][643]=3;
sos_loop[0].somModel.sram_dat[5][644][0]=96'ha4e0;
sos_loop[0].somModel.sram_ptr[5][644]=3;
sos_loop[0].somModel.sram_dat[5][645][0]=96'haede;
sos_loop[0].somModel.sram_ptr[5][645]=3;
sos_loop[0].somModel.sram_dat[5][646][0]=96'hb476;
sos_loop[0].somModel.sram_ptr[5][646]=3;
sos_loop[0].somModel.sram_dat[5][647][0]=96'h4bdf;
sos_loop[0].somModel.sram_ptr[5][647]=3;
sos_loop[0].somModel.sram_dat[5][648][0]=96'h3cb8;
sos_loop[0].somModel.sram_ptr[5][648]=3;
sos_loop[0].somModel.sram_dat[5][649][0]=96'hd010;
sos_loop[0].somModel.sram_ptr[5][649]=3;
sos_loop[0].somModel.sram_dat[5][650][0]=96'h946b;
sos_loop[0].somModel.sram_ptr[5][650]=3;
sos_loop[0].somModel.sram_dat[5][651][0]=96'hafd1;
sos_loop[0].somModel.sram_ptr[5][651]=3;
sos_loop[0].somModel.sram_dat[5][652][0]=96'hf204;
sos_loop[0].somModel.sram_ptr[5][652]=3;
sos_loop[0].somModel.sram_dat[5][653][0]=96'h6781;
sos_loop[0].somModel.sram_ptr[5][653]=3;
sos_loop[0].somModel.sram_dat[5][654][0]=96'hb5f3;
sos_loop[0].somModel.sram_ptr[5][654]=3;
sos_loop[0].somModel.sram_dat[5][655][0]=96'ha278;
sos_loop[0].somModel.sram_ptr[5][655]=3;
sos_loop[0].somModel.sram_dat[5][656][0]=96'h4a51;
sos_loop[0].somModel.sram_ptr[5][656]=3;
sos_loop[0].somModel.sram_dat[5][657][0]=96'hf899;
sos_loop[0].somModel.sram_ptr[5][657]=3;
sos_loop[0].somModel.sram_dat[5][658][0]=96'hed90;
sos_loop[0].somModel.sram_ptr[5][658]=3;
sos_loop[0].somModel.sram_dat[5][659][0]=96'hedf8;
sos_loop[0].somModel.sram_ptr[5][659]=3;
sos_loop[0].somModel.sram_dat[5][660][0]=96'h252e;
sos_loop[0].somModel.sram_ptr[5][660]=3;
sos_loop[0].somModel.sram_dat[5][661][0]=96'h52aa;
sos_loop[0].somModel.sram_ptr[5][661]=3;
sos_loop[0].somModel.sram_dat[5][662][0]=96'h162b;
sos_loop[0].somModel.sram_ptr[5][662]=3;
sos_loop[0].somModel.sram_dat[5][663][0]=96'hfbd9;
sos_loop[0].somModel.sram_ptr[5][663]=3;
sos_loop[0].somModel.sram_dat[5][664][0]=96'h12df;
sos_loop[0].somModel.sram_ptr[5][664]=3;
sos_loop[0].somModel.sram_dat[5][665][0]=96'h7022;
sos_loop[0].somModel.sram_ptr[5][665]=3;
sos_loop[0].somModel.sram_dat[5][666][0]=96'h1a1f;
sos_loop[0].somModel.sram_ptr[5][666]=3;
sos_loop[0].somModel.sram_dat[5][667][0]=96'hf03f;
sos_loop[0].somModel.sram_ptr[5][667]=3;
sos_loop[0].somModel.sram_dat[5][668][0]=96'h324;
sos_loop[0].somModel.sram_ptr[5][668]=3;
sos_loop[0].somModel.sram_dat[5][669][0]=96'h962c;
sos_loop[0].somModel.sram_ptr[5][669]=3;
sos_loop[0].somModel.sram_dat[5][670][0]=96'h3723;
sos_loop[0].somModel.sram_ptr[5][670]=3;
sos_loop[0].somModel.sram_dat[5][671][0]=96'h7c70;
sos_loop[0].somModel.sram_ptr[5][671]=3;
sos_loop[0].somModel.sram_dat[5][672][0]=96'h4bc5;
sos_loop[0].somModel.sram_ptr[5][672]=3;
sos_loop[0].somModel.sram_dat[5][673][0]=96'hca6b;
sos_loop[0].somModel.sram_ptr[5][673]=3;
sos_loop[0].somModel.sram_dat[5][674][0]=96'h6f8b;
sos_loop[0].somModel.sram_ptr[5][674]=3;
sos_loop[0].somModel.sram_dat[5][675][0]=96'h4565;
sos_loop[0].somModel.sram_ptr[5][675]=3;
sos_loop[0].somModel.sram_dat[5][676][0]=96'h3366;
sos_loop[0].somModel.sram_ptr[5][676]=3;
sos_loop[0].somModel.sram_dat[5][677][0]=96'he66a;
sos_loop[0].somModel.sram_ptr[5][677]=3;
sos_loop[0].somModel.sram_dat[5][678][0]=96'h209;
sos_loop[0].somModel.sram_ptr[5][678]=3;
sos_loop[0].somModel.sram_dat[5][679][0]=96'hc785;
sos_loop[0].somModel.sram_ptr[5][679]=3;
sos_loop[0].somModel.sram_dat[5][680][0]=96'hdff4;
sos_loop[0].somModel.sram_ptr[5][680]=3;
sos_loop[0].somModel.sram_dat[5][681][0]=96'h50e;
sos_loop[0].somModel.sram_ptr[5][681]=3;
sos_loop[0].somModel.sram_dat[5][682][0]=96'ha9f5;
sos_loop[0].somModel.sram_ptr[5][682]=3;
sos_loop[0].somModel.sram_dat[5][683][0]=96'hba20;
sos_loop[0].somModel.sram_ptr[5][683]=3;
sos_loop[0].somModel.sram_dat[5][684][0]=96'hba1d;
sos_loop[0].somModel.sram_ptr[5][684]=3;
sos_loop[0].somModel.sram_dat[5][685][0]=96'ha04d;
sos_loop[0].somModel.sram_ptr[5][685]=3;
sos_loop[0].somModel.sram_dat[5][686][0]=96'h5474;
sos_loop[0].somModel.sram_ptr[5][686]=3;
sos_loop[0].somModel.sram_dat[5][687][0]=96'h4961;
sos_loop[0].somModel.sram_ptr[5][687]=3;
sos_loop[0].somModel.sram_dat[5][688][0]=96'hb74e;
sos_loop[0].somModel.sram_ptr[5][688]=3;
sos_loop[0].somModel.sram_dat[5][689][0]=96'he69a;
sos_loop[0].somModel.sram_ptr[5][689]=3;
sos_loop[0].somModel.sram_dat[5][690][0]=96'he108;
sos_loop[0].somModel.sram_ptr[5][690]=3;
sos_loop[0].somModel.sram_dat[5][691][0]=96'h88aa;
sos_loop[0].somModel.sram_ptr[5][691]=3;
sos_loop[0].somModel.sram_dat[5][692][0]=96'hd5b3;
sos_loop[0].somModel.sram_ptr[5][692]=3;
sos_loop[0].somModel.sram_dat[5][693][0]=96'hbb4c;
sos_loop[0].somModel.sram_ptr[5][693]=3;
sos_loop[0].somModel.sram_dat[5][694][0]=96'h9ba6;
sos_loop[0].somModel.sram_ptr[5][694]=3;
sos_loop[0].somModel.sram_dat[5][695][0]=96'h4930;
sos_loop[0].somModel.sram_ptr[5][695]=3;
sos_loop[0].somModel.sram_dat[5][696][0]=96'he153;
sos_loop[0].somModel.sram_ptr[5][696]=3;
sos_loop[0].somModel.sram_dat[5][697][0]=96'h2cbf;
sos_loop[0].somModel.sram_ptr[5][697]=3;
sos_loop[0].somModel.sram_dat[5][698][0]=96'hf52a;
sos_loop[0].somModel.sram_ptr[5][698]=3;
sos_loop[0].somModel.sram_dat[5][699][0]=96'he6da;
sos_loop[0].somModel.sram_ptr[5][699]=3;
sos_loop[0].somModel.sram_dat[5][700][0]=96'he180;
sos_loop[0].somModel.sram_ptr[5][700]=3;
sos_loop[0].somModel.cfg_tbl_sel[5] = 5;
sos_loop[0].somModel.cfg_dat_sel[5] = 4;
sos_loop[0].somModel.cfg_dat_vld[5] = 1;
sos_loop[0].somModel.cfg_miss_ptr[5] = 0;
sos_loop[0].somModel.tcam_data[6][0][0]=80'h00000000000000000000;
sos_loop[0].somModel.tcam_mask[6][0][0]=80'hffffffffffffffffffff;
sos_loop[0].somModel.tcam_data[6][1][0]=80'h00000000c76428a3ac18;
sos_loop[0].somModel.tcam_mask[6][1][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][2][0]=80'h000000006fa2b332a044;
sos_loop[0].somModel.tcam_mask[6][2][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][3][0]=80'h00000000df160ea7e244;
sos_loop[0].somModel.tcam_mask[6][3][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][4][0]=80'h00000000bde8a5158a2b;
sos_loop[0].somModel.tcam_mask[6][4][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][5][0]=80'h000000001c7fcaa5772f;
sos_loop[0].somModel.tcam_mask[6][5][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][6][0]=80'h00000000398bc2065413;
sos_loop[0].somModel.tcam_mask[6][6][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][7][0]=80'h00000000bf26a132d23e;
sos_loop[0].somModel.tcam_mask[6][7][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][8][0]=80'h000000002e5a52ddfb3f;
sos_loop[0].somModel.tcam_mask[6][8][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][9][0]=80'h000000000f9c4f448c4c;
sos_loop[0].somModel.tcam_mask[6][9][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][10][0]=80'h0000000035e4dd182f90;
sos_loop[0].somModel.tcam_mask[6][10][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][11][0]=80'h000000008513d0c50521;
sos_loop[0].somModel.tcam_mask[6][11][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][12][0]=80'h0000000035a66285b62e;
sos_loop[0].somModel.tcam_mask[6][12][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][13][0]=80'h000000004915d9de428f;
sos_loop[0].somModel.tcam_mask[6][13][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][14][0]=80'h000000003eff489073c2;
sos_loop[0].somModel.tcam_mask[6][14][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][15][0]=80'h00000000d00165db49c5;
sos_loop[0].somModel.tcam_mask[6][15][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][16][0]=80'h00000000c6e7d540048a;
sos_loop[0].somModel.tcam_mask[6][16][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][17][0]=80'h000000000d2cf31221e9;
sos_loop[0].somModel.tcam_mask[6][17][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][18][0]=80'h000000009cc2400c08bc;
sos_loop[0].somModel.tcam_mask[6][18][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][19][0]=80'h00000000e84ab68b1a24;
sos_loop[0].somModel.tcam_mask[6][19][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][20][0]=80'h00000000dc9c606e91ae;
sos_loop[0].somModel.tcam_mask[6][20][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][21][0]=80'h000000004b8ee53f7660;
sos_loop[0].somModel.tcam_mask[6][21][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][22][0]=80'h00000000a6dc109cdbbd;
sos_loop[0].somModel.tcam_mask[6][22][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][23][0]=80'h000000002e5acd726cb2;
sos_loop[0].somModel.tcam_mask[6][23][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][24][0]=80'h00000000bb30b2ecd487;
sos_loop[0].somModel.tcam_mask[6][24][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][25][0]=80'h000000009aeec82f8fac;
sos_loop[0].somModel.tcam_mask[6][25][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][26][0]=80'h00000000ab83fe2b985c;
sos_loop[0].somModel.tcam_mask[6][26][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][27][0]=80'h00000000ca3daac02b2f;
sos_loop[0].somModel.tcam_mask[6][27][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][28][0]=80'h000000001a893b2ffa10;
sos_loop[0].somModel.tcam_mask[6][28][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][29][0]=80'h00000000cb1ab883d9ca;
sos_loop[0].somModel.tcam_mask[6][29][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][30][0]=80'h000000006ddb0412e88d;
sos_loop[0].somModel.tcam_mask[6][30][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][31][0]=80'h0000000025d034a677c8;
sos_loop[0].somModel.tcam_mask[6][31][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][32][0]=80'h0000000002ee63ce89af;
sos_loop[0].somModel.tcam_mask[6][32][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[6][33][0]=80'h000000001ab5a710d843;
sos_loop[0].somModel.tcam_mask[6][33][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][34][0]=80'h0000000097e8c062f084;
sos_loop[0].somModel.tcam_mask[6][34][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][35][0]=80'h0000000030a809743d4f;
sos_loop[0].somModel.tcam_mask[6][35][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][36][0]=80'h0000000022420da7f8f4;
sos_loop[0].somModel.tcam_mask[6][36][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][37][0]=80'h00000000afaf284ad3bc;
sos_loop[0].somModel.tcam_mask[6][37][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][38][0]=80'h0000000053bd4f0d7794;
sos_loop[0].somModel.tcam_mask[6][38][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][39][0]=80'h000000005c0d39f2f061;
sos_loop[0].somModel.tcam_mask[6][39][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][40][0]=80'h000000009419a7ce074a;
sos_loop[0].somModel.tcam_mask[6][40][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][41][0]=80'h00000000052d45cc1e4a;
sos_loop[0].somModel.tcam_mask[6][41][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][42][0]=80'h000000009b30665b9971;
sos_loop[0].somModel.tcam_mask[6][42][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][43][0]=80'h0000000020d936f412c1;
sos_loop[0].somModel.tcam_mask[6][43][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][44][0]=80'h000000008b889af41550;
sos_loop[0].somModel.tcam_mask[6][44][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][45][0]=80'h00000000f91ce85e797d;
sos_loop[0].somModel.tcam_mask[6][45][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][46][0]=80'h0000000006e1dbd81191;
sos_loop[0].somModel.tcam_mask[6][46][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][47][0]=80'h00000000345e3c5f1365;
sos_loop[0].somModel.tcam_mask[6][47][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][48][0]=80'h000000008dceefe91dc9;
sos_loop[0].somModel.tcam_mask[6][48][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][49][0]=80'h00000000d47d2191ffed;
sos_loop[0].somModel.tcam_mask[6][49][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][50][0]=80'h000000007d341fbc821b;
sos_loop[0].somModel.tcam_mask[6][50][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][51][0]=80'h000000002e1c5d9ff7d9;
sos_loop[0].somModel.tcam_mask[6][51][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][52][0]=80'h00000000b7c667fd0324;
sos_loop[0].somModel.tcam_mask[6][52][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][53][0]=80'h000000004933bf21a16c;
sos_loop[0].somModel.tcam_mask[6][53][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][54][0]=80'h00000000f9724902347e;
sos_loop[0].somModel.tcam_mask[6][54][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][55][0]=80'h00000000aeb766b220db;
sos_loop[0].somModel.tcam_mask[6][55][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][56][0]=80'h00000000dbbc2a3224ab;
sos_loop[0].somModel.tcam_mask[6][56][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][57][0]=80'h00000000365a679e8085;
sos_loop[0].somModel.tcam_mask[6][57][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][58][0]=80'h00000000eeff7c2b7b33;
sos_loop[0].somModel.tcam_mask[6][58][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][59][0]=80'h0000000045bb6a31bb68;
sos_loop[0].somModel.tcam_mask[6][59][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][60][0]=80'h000000001a81b1c43f91;
sos_loop[0].somModel.tcam_mask[6][60][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][61][0]=80'h000000001de0ad29184a;
sos_loop[0].somModel.tcam_mask[6][61][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][62][0]=80'h000000004eb9229cd415;
sos_loop[0].somModel.tcam_mask[6][62][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][63][0]=80'h0000000075c39cfd15db;
sos_loop[0].somModel.tcam_mask[6][63][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][64][0]=80'h000000000bd7d9ddf726;
sos_loop[0].somModel.tcam_mask[6][64][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][65][0]=80'h00000000788ece7eed43;
sos_loop[0].somModel.tcam_mask[6][65][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][66][0]=80'h00000000689790000fff;
sos_loop[0].somModel.tcam_mask[6][66][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][67][0]=80'h0000000030fca31cf96b;
sos_loop[0].somModel.tcam_mask[6][67][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][68][0]=80'h00000000358975cc2823;
sos_loop[0].somModel.tcam_mask[6][68][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][69][0]=80'h000000006b1cd921c79d;
sos_loop[0].somModel.tcam_mask[6][69][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][70][0]=80'h00000000549a31ff63b7;
sos_loop[0].somModel.tcam_mask[6][70][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][71][0]=80'h00000000310dee607220;
sos_loop[0].somModel.tcam_mask[6][71][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][72][0]=80'h00000000af90fc2fb606;
sos_loop[0].somModel.tcam_mask[6][72][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][73][0]=80'h000000000db655000d3a;
sos_loop[0].somModel.tcam_mask[6][73][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][74][0]=80'h000000008bf35344ab45;
sos_loop[0].somModel.tcam_mask[6][74][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][75][0]=80'h000000002d8a38190b20;
sos_loop[0].somModel.tcam_mask[6][75][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][76][0]=80'h000000000263f7f66582;
sos_loop[0].somModel.tcam_mask[6][76][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[6][77][0]=80'h000000004dfc2ba4768d;
sos_loop[0].somModel.tcam_mask[6][77][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][78][0]=80'h00000000849983bfbe7a;
sos_loop[0].somModel.tcam_mask[6][78][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][79][0]=80'h000000001efcb2f4dd4d;
sos_loop[0].somModel.tcam_mask[6][79][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][80][0]=80'h0000000061e5a9de4569;
sos_loop[0].somModel.tcam_mask[6][80][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][81][0]=80'h00000000770c1c4bd3a5;
sos_loop[0].somModel.tcam_mask[6][81][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][82][0]=80'h00000000500562660aff;
sos_loop[0].somModel.tcam_mask[6][82][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][83][0]=80'h00000000a72a189143e2;
sos_loop[0].somModel.tcam_mask[6][83][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][84][0]=80'h0000000051a64abf0e09;
sos_loop[0].somModel.tcam_mask[6][84][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][85][0]=80'h000000001f5700abe928;
sos_loop[0].somModel.tcam_mask[6][85][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][86][0]=80'h00000000512e72fad6a2;
sos_loop[0].somModel.tcam_mask[6][86][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][87][0]=80'h000000005f3a530396cf;
sos_loop[0].somModel.tcam_mask[6][87][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][88][0]=80'h00000000748487400445;
sos_loop[0].somModel.tcam_mask[6][88][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][89][0]=80'h0000000087719fb3f864;
sos_loop[0].somModel.tcam_mask[6][89][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][90][0]=80'h00000000e88c8f60061d;
sos_loop[0].somModel.tcam_mask[6][90][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][91][0]=80'h000000009f6cc5f93019;
sos_loop[0].somModel.tcam_mask[6][91][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][92][0]=80'h00000000fa9df2c0fa11;
sos_loop[0].somModel.tcam_mask[6][92][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][93][0]=80'h000000003e5de237f4f3;
sos_loop[0].somModel.tcam_mask[6][93][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][94][0]=80'h000000001220e6f8b9fd;
sos_loop[0].somModel.tcam_mask[6][94][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][95][0]=80'h00000000ceb0c2f94c3c;
sos_loop[0].somModel.tcam_mask[6][95][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][96][0]=80'h000000001845b8356ded;
sos_loop[0].somModel.tcam_mask[6][96][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][97][0]=80'h00000000cb7d6f052ed9;
sos_loop[0].somModel.tcam_mask[6][97][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][98][0]=80'h00000000a1d827523dc7;
sos_loop[0].somModel.tcam_mask[6][98][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][99][0]=80'h000000000caf8264a3ea;
sos_loop[0].somModel.tcam_mask[6][99][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][100][0]=80'h0000000038ead3f12916;
sos_loop[0].somModel.tcam_mask[6][100][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][101][0]=80'h0000000013d2ee37c448;
sos_loop[0].somModel.tcam_mask[6][101][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][102][0]=80'h000000003c2fe7d9f34c;
sos_loop[0].somModel.tcam_mask[6][102][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][103][0]=80'h000000003c1db8626079;
sos_loop[0].somModel.tcam_mask[6][103][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][104][0]=80'h00000000865b861ca607;
sos_loop[0].somModel.tcam_mask[6][104][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][105][0]=80'h00000000794600c6d0f4;
sos_loop[0].somModel.tcam_mask[6][105][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][106][0]=80'h00000000e00c57f6e0b3;
sos_loop[0].somModel.tcam_mask[6][106][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][107][0]=80'h00000000e29db65e8903;
sos_loop[0].somModel.tcam_mask[6][107][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][108][0]=80'h000000008e261e6170f3;
sos_loop[0].somModel.tcam_mask[6][108][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][109][0]=80'h0000000066939b10ec73;
sos_loop[0].somModel.tcam_mask[6][109][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][110][0]=80'h0000000070c2e9c3c8eb;
sos_loop[0].somModel.tcam_mask[6][110][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][111][0]=80'h0000000045c66be84cf4;
sos_loop[0].somModel.tcam_mask[6][111][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][112][0]=80'h00000000232cef211d0e;
sos_loop[0].somModel.tcam_mask[6][112][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][113][0]=80'h0000000080542dda5aa2;
sos_loop[0].somModel.tcam_mask[6][113][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][114][0]=80'h00000000474effbc30dd;
sos_loop[0].somModel.tcam_mask[6][114][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][115][0]=80'h00000000e4cebd5c6fa4;
sos_loop[0].somModel.tcam_mask[6][115][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][116][0]=80'h00000000af6a54830375;
sos_loop[0].somModel.tcam_mask[6][116][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][117][0]=80'h000000008ef028be44c1;
sos_loop[0].somModel.tcam_mask[6][117][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][118][0]=80'h000000005fdca8436bf4;
sos_loop[0].somModel.tcam_mask[6][118][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][119][0]=80'h000000006e7e1c15bd08;
sos_loop[0].somModel.tcam_mask[6][119][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][120][0]=80'h00000000134c1f65fd66;
sos_loop[0].somModel.tcam_mask[6][120][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][121][0]=80'h00000000cea87493679f;
sos_loop[0].somModel.tcam_mask[6][121][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][122][0]=80'h00000000ceb7bc309c1a;
sos_loop[0].somModel.tcam_mask[6][122][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][123][0]=80'h0000000061a6f8771878;
sos_loop[0].somModel.tcam_mask[6][123][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][124][0]=80'h00000000cedef6a567fe;
sos_loop[0].somModel.tcam_mask[6][124][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][125][0]=80'h000000002e32a08622cd;
sos_loop[0].somModel.tcam_mask[6][125][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][126][0]=80'h000000005356e16b8fd7;
sos_loop[0].somModel.tcam_mask[6][126][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][127][0]=80'h00000000fd605bd942c3;
sos_loop[0].somModel.tcam_mask[6][127][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][128][0]=80'h0000000000d5f103f449;
sos_loop[0].somModel.tcam_mask[6][128][0]=80'hffffffffff0000000000;
sos_loop[0].somModel.tcam_data[6][129][0]=80'h000000005f57f4362b22;
sos_loop[0].somModel.tcam_mask[6][129][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][130][0]=80'h000000002e67f284f871;
sos_loop[0].somModel.tcam_mask[6][130][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][131][0]=80'h00000000ecd79dcadc01;
sos_loop[0].somModel.tcam_mask[6][131][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][132][0]=80'h00000000e00525c7b0f8;
sos_loop[0].somModel.tcam_mask[6][132][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][133][0]=80'h00000000b3cf483e6c80;
sos_loop[0].somModel.tcam_mask[6][133][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][134][0]=80'h0000000077eb26f31bbe;
sos_loop[0].somModel.tcam_mask[6][134][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][135][0]=80'h000000008b676c49d915;
sos_loop[0].somModel.tcam_mask[6][135][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][136][0]=80'h000000000a2822acbd35;
sos_loop[0].somModel.tcam_mask[6][136][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][137][0]=80'h0000000003a257929df1;
sos_loop[0].somModel.tcam_mask[6][137][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[6][138][0]=80'h00000000e9b0e1c40a18;
sos_loop[0].somModel.tcam_mask[6][138][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][139][0]=80'h000000003f10a0b32f42;
sos_loop[0].somModel.tcam_mask[6][139][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][140][0]=80'h00000000f8a042a8b1d1;
sos_loop[0].somModel.tcam_mask[6][140][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][141][0]=80'h00000000c010041f98fe;
sos_loop[0].somModel.tcam_mask[6][141][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][142][0]=80'h000000006f5155d6bf2a;
sos_loop[0].somModel.tcam_mask[6][142][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][143][0]=80'h000000006174e0aee88e;
sos_loop[0].somModel.tcam_mask[6][143][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][144][0]=80'h00000000d8f296505931;
sos_loop[0].somModel.tcam_mask[6][144][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][145][0]=80'h00000000e512e3c64789;
sos_loop[0].somModel.tcam_mask[6][145][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][146][0]=80'h00000000373e0b9976b9;
sos_loop[0].somModel.tcam_mask[6][146][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][147][0]=80'h0000000003e7dacda18b;
sos_loop[0].somModel.tcam_mask[6][147][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[6][148][0]=80'h000000000964ddbc00a5;
sos_loop[0].somModel.tcam_mask[6][148][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][149][0]=80'h0000000054781b947c65;
sos_loop[0].somModel.tcam_mask[6][149][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][150][0]=80'h000000004e476ae23070;
sos_loop[0].somModel.tcam_mask[6][150][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][151][0]=80'h00000000965a202c5dd1;
sos_loop[0].somModel.tcam_mask[6][151][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][152][0]=80'h000000006eeef25e5a0e;
sos_loop[0].somModel.tcam_mask[6][152][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][153][0]=80'h00000000bd9be825e53c;
sos_loop[0].somModel.tcam_mask[6][153][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][154][0]=80'h000000005a0d2b0e2652;
sos_loop[0].somModel.tcam_mask[6][154][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][155][0]=80'h00000000f02c2960a78f;
sos_loop[0].somModel.tcam_mask[6][155][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][156][0]=80'h0000000043801573ed5c;
sos_loop[0].somModel.tcam_mask[6][156][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][157][0]=80'h0000000034d1a3628645;
sos_loop[0].somModel.tcam_mask[6][157][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][158][0]=80'h00000000476d2c7ebc16;
sos_loop[0].somModel.tcam_mask[6][158][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][159][0]=80'h00000000a17de6c9b9c6;
sos_loop[0].somModel.tcam_mask[6][159][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][160][0]=80'h000000002e3b2da7cb0e;
sos_loop[0].somModel.tcam_mask[6][160][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][161][0]=80'h00000000618fe75b3a00;
sos_loop[0].somModel.tcam_mask[6][161][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][162][0]=80'h000000007868e9b929a2;
sos_loop[0].somModel.tcam_mask[6][162][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][163][0]=80'h00000000cbe5e4137d1a;
sos_loop[0].somModel.tcam_mask[6][163][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][164][0]=80'h000000006771e8c490b5;
sos_loop[0].somModel.tcam_mask[6][164][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][165][0]=80'h000000007be9cc15dbad;
sos_loop[0].somModel.tcam_mask[6][165][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][166][0]=80'h000000008c89b097b14c;
sos_loop[0].somModel.tcam_mask[6][166][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][167][0]=80'h00000000f2124342ae18;
sos_loop[0].somModel.tcam_mask[6][167][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][168][0]=80'h00000000330261ba3670;
sos_loop[0].somModel.tcam_mask[6][168][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][169][0]=80'h0000000042c4edb6d896;
sos_loop[0].somModel.tcam_mask[6][169][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][170][0]=80'h0000000023a570bc32da;
sos_loop[0].somModel.tcam_mask[6][170][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][171][0]=80'h00000000db4f2973fc73;
sos_loop[0].somModel.tcam_mask[6][171][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][172][0]=80'h000000004c40d88318b1;
sos_loop[0].somModel.tcam_mask[6][172][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][173][0]=80'h000000001273739101e3;
sos_loop[0].somModel.tcam_mask[6][173][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][174][0]=80'h000000009c2ebac8770d;
sos_loop[0].somModel.tcam_mask[6][174][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][175][0]=80'h00000000aaeaffde1744;
sos_loop[0].somModel.tcam_mask[6][175][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][176][0]=80'h0000000067b1d0406ac4;
sos_loop[0].somModel.tcam_mask[6][176][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][177][0]=80'h00000000602be7c25423;
sos_loop[0].somModel.tcam_mask[6][177][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][178][0]=80'h000000007bd2374d89da;
sos_loop[0].somModel.tcam_mask[6][178][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][179][0]=80'h00000000484efbf68ee5;
sos_loop[0].somModel.tcam_mask[6][179][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][180][0]=80'h000000008c2970d5df55;
sos_loop[0].somModel.tcam_mask[6][180][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][181][0]=80'h00000000aec65cebfe7b;
sos_loop[0].somModel.tcam_mask[6][181][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][182][0]=80'h0000000094dfc4cad63a;
sos_loop[0].somModel.tcam_mask[6][182][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][183][0]=80'h0000000016398c9c5329;
sos_loop[0].somModel.tcam_mask[6][183][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][184][0]=80'h00000000c1d9c5b84501;
sos_loop[0].somModel.tcam_mask[6][184][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][185][0]=80'h00000000d1ad3332662b;
sos_loop[0].somModel.tcam_mask[6][185][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][186][0]=80'h00000000b91d094ca5fa;
sos_loop[0].somModel.tcam_mask[6][186][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][187][0]=80'h0000000066807169ce5b;
sos_loop[0].somModel.tcam_mask[6][187][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][188][0]=80'h000000006ef096e4f564;
sos_loop[0].somModel.tcam_mask[6][188][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][189][0]=80'h00000000328864e675f7;
sos_loop[0].somModel.tcam_mask[6][189][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][190][0]=80'h000000007dae2b0e1b45;
sos_loop[0].somModel.tcam_mask[6][190][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][191][0]=80'h00000000bcb94b47b6e1;
sos_loop[0].somModel.tcam_mask[6][191][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][192][0]=80'h00000000969630df4be5;
sos_loop[0].somModel.tcam_mask[6][192][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][193][0]=80'h000000008fa1021a531a;
sos_loop[0].somModel.tcam_mask[6][193][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][194][0]=80'h00000000872d61d5debf;
sos_loop[0].somModel.tcam_mask[6][194][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][195][0]=80'h00000000991610788933;
sos_loop[0].somModel.tcam_mask[6][195][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][196][0]=80'h000000000abf899e0a35;
sos_loop[0].somModel.tcam_mask[6][196][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][197][0]=80'h000000009a50b37b4c4e;
sos_loop[0].somModel.tcam_mask[6][197][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][198][0]=80'h00000000a57859f9c477;
sos_loop[0].somModel.tcam_mask[6][198][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][199][0]=80'h000000000079cd60c49c;
sos_loop[0].somModel.tcam_mask[6][199][0]=80'hffffffffff8000000000;
sos_loop[0].somModel.tcam_data[6][200][0]=80'h00000000116a5a1abd7d;
sos_loop[0].somModel.tcam_mask[6][200][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][201][0]=80'h00000000c21fd0b46818;
sos_loop[0].somModel.tcam_mask[6][201][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][202][0]=80'h00000000cb7c1d8cfffa;
sos_loop[0].somModel.tcam_mask[6][202][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][203][0]=80'h000000005da2668e789f;
sos_loop[0].somModel.tcam_mask[6][203][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][204][0]=80'h00000000a975554d1660;
sos_loop[0].somModel.tcam_mask[6][204][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][205][0]=80'h00000000f527f8412a24;
sos_loop[0].somModel.tcam_mask[6][205][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][206][0]=80'h000000006e7cabe12a47;
sos_loop[0].somModel.tcam_mask[6][206][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][207][0]=80'h00000000ecce1c4cd86e;
sos_loop[0].somModel.tcam_mask[6][207][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][208][0]=80'h0000000072d3d3fcd72b;
sos_loop[0].somModel.tcam_mask[6][208][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][209][0]=80'h00000000839e1fb55d44;
sos_loop[0].somModel.tcam_mask[6][209][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][210][0]=80'h00000000478398e0b9ee;
sos_loop[0].somModel.tcam_mask[6][210][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][211][0]=80'h000000008530d50e759f;
sos_loop[0].somModel.tcam_mask[6][211][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][212][0]=80'h0000000011f968361ebd;
sos_loop[0].somModel.tcam_mask[6][212][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][213][0]=80'h000000008ce994cc083f;
sos_loop[0].somModel.tcam_mask[6][213][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][214][0]=80'h000000002c23f84988ee;
sos_loop[0].somModel.tcam_mask[6][214][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][215][0]=80'h000000009760938f25c2;
sos_loop[0].somModel.tcam_mask[6][215][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][216][0]=80'h00000000274efbfa8211;
sos_loop[0].somModel.tcam_mask[6][216][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][217][0]=80'h00000000694132b93ba3;
sos_loop[0].somModel.tcam_mask[6][217][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][218][0]=80'h000000000682f3056401;
sos_loop[0].somModel.tcam_mask[6][218][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][219][0]=80'h00000000d1c36a785d4f;
sos_loop[0].somModel.tcam_mask[6][219][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][220][0]=80'h000000004ae9b6d2ef4f;
sos_loop[0].somModel.tcam_mask[6][220][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][221][0]=80'h00000000c9c32ab41eeb;
sos_loop[0].somModel.tcam_mask[6][221][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][222][0]=80'h00000000cbc076ebe28e;
sos_loop[0].somModel.tcam_mask[6][222][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][223][0]=80'h00000000fbda31fd76c0;
sos_loop[0].somModel.tcam_mask[6][223][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][224][0]=80'h000000009a099a151b35;
sos_loop[0].somModel.tcam_mask[6][224][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][225][0]=80'h0000000054a1681b3ffb;
sos_loop[0].somModel.tcam_mask[6][225][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][226][0]=80'h00000000f0cf8f9ee272;
sos_loop[0].somModel.tcam_mask[6][226][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][227][0]=80'h000000003f535b44d28a;
sos_loop[0].somModel.tcam_mask[6][227][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][228][0]=80'h000000007ae44fa333c8;
sos_loop[0].somModel.tcam_mask[6][228][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][229][0]=80'h00000000b665ce7f735a;
sos_loop[0].somModel.tcam_mask[6][229][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][230][0]=80'h00000000626c7ae8774d;
sos_loop[0].somModel.tcam_mask[6][230][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][231][0]=80'h00000000f3cddb51d392;
sos_loop[0].somModel.tcam_mask[6][231][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][232][0]=80'h00000000944a75a8319c;
sos_loop[0].somModel.tcam_mask[6][232][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][233][0]=80'h00000000eaacb9890fae;
sos_loop[0].somModel.tcam_mask[6][233][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][234][0]=80'h00000000046f6540ec7f;
sos_loop[0].somModel.tcam_mask[6][234][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][235][0]=80'h00000000c6088fc1bd3d;
sos_loop[0].somModel.tcam_mask[6][235][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][236][0]=80'h000000005e0b61c56031;
sos_loop[0].somModel.tcam_mask[6][236][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][237][0]=80'h00000000027b4c51c3bb;
sos_loop[0].somModel.tcam_mask[6][237][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[6][238][0]=80'h00000000be4d82d7e60e;
sos_loop[0].somModel.tcam_mask[6][238][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][239][0]=80'h000000007eef6a0932c5;
sos_loop[0].somModel.tcam_mask[6][239][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][240][0]=80'h00000000564f40cb3bc6;
sos_loop[0].somModel.tcam_mask[6][240][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][241][0]=80'h0000000049ba0e14ede1;
sos_loop[0].somModel.tcam_mask[6][241][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][242][0]=80'h000000000ffa1385e8e1;
sos_loop[0].somModel.tcam_mask[6][242][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][243][0]=80'h00000000c2a6a6c5875c;
sos_loop[0].somModel.tcam_mask[6][243][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][244][0]=80'h0000000046ed88992ff9;
sos_loop[0].somModel.tcam_mask[6][244][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][245][0]=80'h000000007bd52c488741;
sos_loop[0].somModel.tcam_mask[6][245][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][246][0]=80'h00000000dd037b320186;
sos_loop[0].somModel.tcam_mask[6][246][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][247][0]=80'h00000000bc45bae8ac0a;
sos_loop[0].somModel.tcam_mask[6][247][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][248][0]=80'h000000005b06c7e96f30;
sos_loop[0].somModel.tcam_mask[6][248][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][249][0]=80'h00000000d4ddc557a673;
sos_loop[0].somModel.tcam_mask[6][249][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][250][0]=80'h0000000053ec21af6aa7;
sos_loop[0].somModel.tcam_mask[6][250][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][251][0]=80'h0000000017ac57f88e87;
sos_loop[0].somModel.tcam_mask[6][251][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][252][0]=80'h00000000a4100e4032cc;
sos_loop[0].somModel.tcam_mask[6][252][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][253][0]=80'h00000000140fa51dda60;
sos_loop[0].somModel.tcam_mask[6][253][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][254][0]=80'h00000000ba76b63b04af;
sos_loop[0].somModel.tcam_mask[6][254][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][255][0]=80'h000000007bf30212d42d;
sos_loop[0].somModel.tcam_mask[6][255][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][256][0]=80'h00000000389a856d0929;
sos_loop[0].somModel.tcam_mask[6][256][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][257][0]=80'h00000000971def77bfa0;
sos_loop[0].somModel.tcam_mask[6][257][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][258][0]=80'h000000007fea6ca2dda9;
sos_loop[0].somModel.tcam_mask[6][258][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][259][0]=80'h000000006cc87b7163e1;
sos_loop[0].somModel.tcam_mask[6][259][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][260][0]=80'h00000000652f37432033;
sos_loop[0].somModel.tcam_mask[6][260][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][261][0]=80'h0000000094ca0afeaf40;
sos_loop[0].somModel.tcam_mask[6][261][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][262][0]=80'h00000000aa6075a82cfd;
sos_loop[0].somModel.tcam_mask[6][262][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][263][0]=80'h00000000e393132fbd4d;
sos_loop[0].somModel.tcam_mask[6][263][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][264][0]=80'h000000008617fb8769a3;
sos_loop[0].somModel.tcam_mask[6][264][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][265][0]=80'h00000000d45704f554fa;
sos_loop[0].somModel.tcam_mask[6][265][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][266][0]=80'h00000000083aeac67707;
sos_loop[0].somModel.tcam_mask[6][266][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][267][0]=80'h00000000ad11dd592c9a;
sos_loop[0].somModel.tcam_mask[6][267][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][268][0]=80'h00000000199fcd09ed28;
sos_loop[0].somModel.tcam_mask[6][268][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][269][0]=80'h00000000306fc67d4fd2;
sos_loop[0].somModel.tcam_mask[6][269][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][270][0]=80'h00000000ded308236673;
sos_loop[0].somModel.tcam_mask[6][270][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][271][0]=80'h000000006bb4f3981543;
sos_loop[0].somModel.tcam_mask[6][271][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][272][0]=80'h0000000028d774fa8bab;
sos_loop[0].somModel.tcam_mask[6][272][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][273][0]=80'h000000005f39e126fa40;
sos_loop[0].somModel.tcam_mask[6][273][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][274][0]=80'h000000004ec1930dd830;
sos_loop[0].somModel.tcam_mask[6][274][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][275][0]=80'h000000002eabafa47444;
sos_loop[0].somModel.tcam_mask[6][275][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][276][0]=80'h00000000f2c4354979b5;
sos_loop[0].somModel.tcam_mask[6][276][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][277][0]=80'h000000004375ff2839ff;
sos_loop[0].somModel.tcam_mask[6][277][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][278][0]=80'h00000000831847d750e3;
sos_loop[0].somModel.tcam_mask[6][278][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][279][0]=80'h000000006d4ff70a7fc3;
sos_loop[0].somModel.tcam_mask[6][279][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][280][0]=80'h0000000067633ad96690;
sos_loop[0].somModel.tcam_mask[6][280][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][281][0]=80'h0000000058b1bb7ab35b;
sos_loop[0].somModel.tcam_mask[6][281][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][282][0]=80'h00000000378d65b1297a;
sos_loop[0].somModel.tcam_mask[6][282][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][283][0]=80'h000000008ab24a720a34;
sos_loop[0].somModel.tcam_mask[6][283][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][284][0]=80'h000000009b617faf808a;
sos_loop[0].somModel.tcam_mask[6][284][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][285][0]=80'h000000002b5be33345f9;
sos_loop[0].somModel.tcam_mask[6][285][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][286][0]=80'h0000000080b069925240;
sos_loop[0].somModel.tcam_mask[6][286][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][287][0]=80'h0000000064819ae5ce38;
sos_loop[0].somModel.tcam_mask[6][287][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][288][0]=80'h00000000c8a2886319ad;
sos_loop[0].somModel.tcam_mask[6][288][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][289][0]=80'h00000000bba80680cd74;
sos_loop[0].somModel.tcam_mask[6][289][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][290][0]=80'h00000000c624c1780420;
sos_loop[0].somModel.tcam_mask[6][290][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][291][0]=80'h000000000df4dc19f8a0;
sos_loop[0].somModel.tcam_mask[6][291][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][292][0]=80'h00000000bf4fc4c5109d;
sos_loop[0].somModel.tcam_mask[6][292][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][293][0]=80'h00000000230e53a6e40d;
sos_loop[0].somModel.tcam_mask[6][293][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][294][0]=80'h000000006a8845704812;
sos_loop[0].somModel.tcam_mask[6][294][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][295][0]=80'h00000000d02d7e61c3ff;
sos_loop[0].somModel.tcam_mask[6][295][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][296][0]=80'h0000000042d9ad4b7cb5;
sos_loop[0].somModel.tcam_mask[6][296][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][297][0]=80'h000000006620c43e40cd;
sos_loop[0].somModel.tcam_mask[6][297][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][298][0]=80'h00000000572b2a5075a9;
sos_loop[0].somModel.tcam_mask[6][298][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][299][0]=80'h000000000bc0a3cd8632;
sos_loop[0].somModel.tcam_mask[6][299][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][300][0]=80'h00000000318840f45c23;
sos_loop[0].somModel.tcam_mask[6][300][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][301][0]=80'h000000007ec0b9f2df84;
sos_loop[0].somModel.tcam_mask[6][301][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][302][0]=80'h000000000708eaeea371;
sos_loop[0].somModel.tcam_mask[6][302][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][303][0]=80'h0000000029e3e9901c1f;
sos_loop[0].somModel.tcam_mask[6][303][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][304][0]=80'h00000000f4f0fb40376f;
sos_loop[0].somModel.tcam_mask[6][304][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][305][0]=80'h000000007de8c27c7bf8;
sos_loop[0].somModel.tcam_mask[6][305][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][306][0]=80'h00000000722214538bb3;
sos_loop[0].somModel.tcam_mask[6][306][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][307][0]=80'h00000000b35284a2e8f3;
sos_loop[0].somModel.tcam_mask[6][307][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][308][0]=80'h00000000c1e963dc4088;
sos_loop[0].somModel.tcam_mask[6][308][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][309][0]=80'h0000000050d5503770e6;
sos_loop[0].somModel.tcam_mask[6][309][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][310][0]=80'h00000000b63951662a30;
sos_loop[0].somModel.tcam_mask[6][310][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][311][0]=80'h000000007eddea567619;
sos_loop[0].somModel.tcam_mask[6][311][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][312][0]=80'h000000004eab0a109e8f;
sos_loop[0].somModel.tcam_mask[6][312][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][313][0]=80'h00000000e549f26a551a;
sos_loop[0].somModel.tcam_mask[6][313][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][314][0]=80'h00000000161e12d7d5f4;
sos_loop[0].somModel.tcam_mask[6][314][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][315][0]=80'h000000002fb8691cf03d;
sos_loop[0].somModel.tcam_mask[6][315][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][316][0]=80'h000000006d0dd414bd88;
sos_loop[0].somModel.tcam_mask[6][316][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][317][0]=80'h00000000d47f0cfd8269;
sos_loop[0].somModel.tcam_mask[6][317][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][318][0]=80'h00000000e7fe58f76aac;
sos_loop[0].somModel.tcam_mask[6][318][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][319][0]=80'h00000000cddb5437e4b9;
sos_loop[0].somModel.tcam_mask[6][319][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][320][0]=80'h0000000058ac2d7d65c1;
sos_loop[0].somModel.tcam_mask[6][320][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][321][0]=80'h00000000e81d8eb85034;
sos_loop[0].somModel.tcam_mask[6][321][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][322][0]=80'h00000000a6fb99d69d1b;
sos_loop[0].somModel.tcam_mask[6][322][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][323][0]=80'h0000000085db0f2ad52e;
sos_loop[0].somModel.tcam_mask[6][323][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][324][0]=80'h00000000ba447f49c0b1;
sos_loop[0].somModel.tcam_mask[6][324][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][325][0]=80'h0000000099d3496acd35;
sos_loop[0].somModel.tcam_mask[6][325][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][326][0]=80'h0000000040e7e1b07303;
sos_loop[0].somModel.tcam_mask[6][326][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][327][0]=80'h0000000055f948ebe91d;
sos_loop[0].somModel.tcam_mask[6][327][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][328][0]=80'h00000000392c0459ce02;
sos_loop[0].somModel.tcam_mask[6][328][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][329][0]=80'h000000007e3d419f5d34;
sos_loop[0].somModel.tcam_mask[6][329][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][330][0]=80'h00000000e74efb58eaa7;
sos_loop[0].somModel.tcam_mask[6][330][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][331][0]=80'h00000000f83f581e4482;
sos_loop[0].somModel.tcam_mask[6][331][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][332][0]=80'h000000009cce1dfeef14;
sos_loop[0].somModel.tcam_mask[6][332][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][333][0]=80'h000000004b70936e9f64;
sos_loop[0].somModel.tcam_mask[6][333][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][334][0]=80'h000000008f60bf446783;
sos_loop[0].somModel.tcam_mask[6][334][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][335][0]=80'h0000000093a9046448e2;
sos_loop[0].somModel.tcam_mask[6][335][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][336][0]=80'h000000006e3ce4ac6730;
sos_loop[0].somModel.tcam_mask[6][336][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][337][0]=80'h0000000084de22fbc40a;
sos_loop[0].somModel.tcam_mask[6][337][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][338][0]=80'h000000002d98732c0914;
sos_loop[0].somModel.tcam_mask[6][338][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][339][0]=80'h00000000588e0584287c;
sos_loop[0].somModel.tcam_mask[6][339][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][340][0]=80'h000000008f50e0497e89;
sos_loop[0].somModel.tcam_mask[6][340][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][341][0]=80'h00000000b0e119fb2555;
sos_loop[0].somModel.tcam_mask[6][341][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][342][0]=80'h000000004cd3c2cde21a;
sos_loop[0].somModel.tcam_mask[6][342][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][343][0]=80'h00000000da342cb3beee;
sos_loop[0].somModel.tcam_mask[6][343][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][344][0]=80'h000000009f7fc5e6a042;
sos_loop[0].somModel.tcam_mask[6][344][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][345][0]=80'h00000000cc5300c82669;
sos_loop[0].somModel.tcam_mask[6][345][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][346][0]=80'h000000006a1ec386bf00;
sos_loop[0].somModel.tcam_mask[6][346][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][347][0]=80'h000000002317e8d90545;
sos_loop[0].somModel.tcam_mask[6][347][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][348][0]=80'h000000008d4fe98625cf;
sos_loop[0].somModel.tcam_mask[6][348][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][349][0]=80'h00000000060665e2c19e;
sos_loop[0].somModel.tcam_mask[6][349][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][350][0]=80'h00000000596674fbbfb1;
sos_loop[0].somModel.tcam_mask[6][350][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][351][0]=80'h000000005c7688d8aad5;
sos_loop[0].somModel.tcam_mask[6][351][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][352][0]=80'h0000000099c3cb202d30;
sos_loop[0].somModel.tcam_mask[6][352][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][353][0]=80'h00000000a86ac83a7681;
sos_loop[0].somModel.tcam_mask[6][353][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][354][0]=80'h00000000f9f330aaf7e5;
sos_loop[0].somModel.tcam_mask[6][354][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][355][0]=80'h000000003c3dcdb988e5;
sos_loop[0].somModel.tcam_mask[6][355][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][356][0]=80'h0000000082440e73e0a4;
sos_loop[0].somModel.tcam_mask[6][356][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][357][0]=80'h00000000deb63d376bdd;
sos_loop[0].somModel.tcam_mask[6][357][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][358][0]=80'h000000003f13c6d986da;
sos_loop[0].somModel.tcam_mask[6][358][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][359][0]=80'h00000000959a11161a8a;
sos_loop[0].somModel.tcam_mask[6][359][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][360][0]=80'h0000000004fc4b9709a2;
sos_loop[0].somModel.tcam_mask[6][360][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][361][0]=80'h000000000603260a4fa8;
sos_loop[0].somModel.tcam_mask[6][361][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][362][0]=80'h00000000317642426d30;
sos_loop[0].somModel.tcam_mask[6][362][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][363][0]=80'h0000000093eea5159da0;
sos_loop[0].somModel.tcam_mask[6][363][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][364][0]=80'h00000000a6a6c5effbb8;
sos_loop[0].somModel.tcam_mask[6][364][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][365][0]=80'h000000009a556fc0f1e1;
sos_loop[0].somModel.tcam_mask[6][365][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][366][0]=80'h00000000ca8bfde422b1;
sos_loop[0].somModel.tcam_mask[6][366][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][367][0]=80'h000000006b3d4da4a0e4;
sos_loop[0].somModel.tcam_mask[6][367][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][368][0]=80'h00000000b8725432eee0;
sos_loop[0].somModel.tcam_mask[6][368][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][369][0]=80'h000000002a5f4d97572c;
sos_loop[0].somModel.tcam_mask[6][369][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][370][0]=80'h0000000003f4b2f37c91;
sos_loop[0].somModel.tcam_mask[6][370][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[6][371][0]=80'h000000006d012a56f306;
sos_loop[0].somModel.tcam_mask[6][371][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][372][0]=80'h00000000f39c18ff7423;
sos_loop[0].somModel.tcam_mask[6][372][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][373][0]=80'h0000000064fe54c3d020;
sos_loop[0].somModel.tcam_mask[6][373][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][374][0]=80'h000000005941386df853;
sos_loop[0].somModel.tcam_mask[6][374][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][375][0]=80'h00000000fd5081a7023d;
sos_loop[0].somModel.tcam_mask[6][375][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][376][0]=80'h0000000059d252677e44;
sos_loop[0].somModel.tcam_mask[6][376][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][377][0]=80'h00000000b1ef710456c8;
sos_loop[0].somModel.tcam_mask[6][377][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][378][0]=80'h000000008a3b29afa55f;
sos_loop[0].somModel.tcam_mask[6][378][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][379][0]=80'h00000000a8f4af7c920a;
sos_loop[0].somModel.tcam_mask[6][379][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][380][0]=80'h000000009b5b556528f0;
sos_loop[0].somModel.tcam_mask[6][380][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][381][0]=80'h000000008d75c4ce6384;
sos_loop[0].somModel.tcam_mask[6][381][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][382][0]=80'h00000000644e172a4d39;
sos_loop[0].somModel.tcam_mask[6][382][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][383][0]=80'h000000004e2c31c4e9bf;
sos_loop[0].somModel.tcam_mask[6][383][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][384][0]=80'h00000000fb16e104670e;
sos_loop[0].somModel.tcam_mask[6][384][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][385][0]=80'h00000000edda66338267;
sos_loop[0].somModel.tcam_mask[6][385][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][386][0]=80'h00000000028c12a16f1b;
sos_loop[0].somModel.tcam_mask[6][386][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[6][387][0]=80'h00000000ff84824ad314;
sos_loop[0].somModel.tcam_mask[6][387][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][388][0]=80'h000000000be7756aeeab;
sos_loop[0].somModel.tcam_mask[6][388][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][389][0]=80'h000000007e61e055303f;
sos_loop[0].somModel.tcam_mask[6][389][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][390][0]=80'h00000000aac7193a22af;
sos_loop[0].somModel.tcam_mask[6][390][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][391][0]=80'h00000000565f0106873e;
sos_loop[0].somModel.tcam_mask[6][391][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][392][0]=80'h0000000075032e61802d;
sos_loop[0].somModel.tcam_mask[6][392][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][393][0]=80'h00000000f2f7c9dbbf6e;
sos_loop[0].somModel.tcam_mask[6][393][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][394][0]=80'h00000000c616b82074dc;
sos_loop[0].somModel.tcam_mask[6][394][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][395][0]=80'h000000009b90c73a26b9;
sos_loop[0].somModel.tcam_mask[6][395][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][396][0]=80'h00000000f1aad48501e0;
sos_loop[0].somModel.tcam_mask[6][396][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][397][0]=80'h00000000b50e5a5b2331;
sos_loop[0].somModel.tcam_mask[6][397][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][398][0]=80'h000000000536e70ff511;
sos_loop[0].somModel.tcam_mask[6][398][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][399][0]=80'h00000000500f137223d6;
sos_loop[0].somModel.tcam_mask[6][399][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][400][0]=80'h000000002791051b62a6;
sos_loop[0].somModel.tcam_mask[6][400][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][401][0]=80'h00000000c4eb2c045df0;
sos_loop[0].somModel.tcam_mask[6][401][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][402][0]=80'h00000000a4ad1b4e4c65;
sos_loop[0].somModel.tcam_mask[6][402][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][403][0]=80'h000000005dcd203c62ab;
sos_loop[0].somModel.tcam_mask[6][403][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][404][0]=80'h00000000bd2053fe1aa1;
sos_loop[0].somModel.tcam_mask[6][404][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][405][0]=80'h00000000dd873733eebd;
sos_loop[0].somModel.tcam_mask[6][405][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][406][0]=80'h00000000d5cc8944cc44;
sos_loop[0].somModel.tcam_mask[6][406][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][407][0]=80'h00000000df75e34c1d60;
sos_loop[0].somModel.tcam_mask[6][407][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][408][0]=80'h0000000069516c90e02b;
sos_loop[0].somModel.tcam_mask[6][408][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][409][0]=80'h00000000ba7434218648;
sos_loop[0].somModel.tcam_mask[6][409][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][410][0]=80'h0000000075995e082cc9;
sos_loop[0].somModel.tcam_mask[6][410][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][411][0]=80'h000000008f8a0618c492;
sos_loop[0].somModel.tcam_mask[6][411][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][412][0]=80'h0000000085652adefb50;
sos_loop[0].somModel.tcam_mask[6][412][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][413][0]=80'h0000000084e3bbb346a9;
sos_loop[0].somModel.tcam_mask[6][413][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][414][0]=80'h00000000ce288545ff5c;
sos_loop[0].somModel.tcam_mask[6][414][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][415][0]=80'h00000000f34840529bc7;
sos_loop[0].somModel.tcam_mask[6][415][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][416][0]=80'h0000000093b680734ca8;
sos_loop[0].somModel.tcam_mask[6][416][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][417][0]=80'h000000006d3e5930bf31;
sos_loop[0].somModel.tcam_mask[6][417][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][418][0]=80'h000000004c6bb4e13dd2;
sos_loop[0].somModel.tcam_mask[6][418][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][419][0]=80'h00000000c17e7cae146d;
sos_loop[0].somModel.tcam_mask[6][419][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][420][0]=80'h000000003a01e234f448;
sos_loop[0].somModel.tcam_mask[6][420][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][421][0]=80'h000000001f6089a70d31;
sos_loop[0].somModel.tcam_mask[6][421][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][422][0]=80'h00000000e9910acedf01;
sos_loop[0].somModel.tcam_mask[6][422][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][423][0]=80'h0000000092c1be63a45c;
sos_loop[0].somModel.tcam_mask[6][423][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][424][0]=80'h0000000077250b5545e8;
sos_loop[0].somModel.tcam_mask[6][424][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][425][0]=80'h0000000041875a4af1b4;
sos_loop[0].somModel.tcam_mask[6][425][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][426][0]=80'h000000001f7188b8f195;
sos_loop[0].somModel.tcam_mask[6][426][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][427][0]=80'h00000000e7043697f5e9;
sos_loop[0].somModel.tcam_mask[6][427][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][428][0]=80'h00000000ccb0a5325cbe;
sos_loop[0].somModel.tcam_mask[6][428][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][429][0]=80'h00000000f77c99d0ae10;
sos_loop[0].somModel.tcam_mask[6][429][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][430][0]=80'h0000000051c66267cec7;
sos_loop[0].somModel.tcam_mask[6][430][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][431][0]=80'h00000000a3eb7b517f7d;
sos_loop[0].somModel.tcam_mask[6][431][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][432][0]=80'h000000005e4b84a9a324;
sos_loop[0].somModel.tcam_mask[6][432][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][433][0]=80'h00000000263366d9a934;
sos_loop[0].somModel.tcam_mask[6][433][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][434][0]=80'h0000000035cd167e2bad;
sos_loop[0].somModel.tcam_mask[6][434][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][435][0]=80'h000000000b2c3bbf8fba;
sos_loop[0].somModel.tcam_mask[6][435][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][436][0]=80'h000000008f19a66976c7;
sos_loop[0].somModel.tcam_mask[6][436][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][437][0]=80'h00000000e0b42c35622b;
sos_loop[0].somModel.tcam_mask[6][437][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][438][0]=80'h00000000dca9a6f1782c;
sos_loop[0].somModel.tcam_mask[6][438][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][439][0]=80'h000000009a1541c274a2;
sos_loop[0].somModel.tcam_mask[6][439][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][440][0]=80'h0000000044768a38b95d;
sos_loop[0].somModel.tcam_mask[6][440][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][441][0]=80'h0000000038f48a68b142;
sos_loop[0].somModel.tcam_mask[6][441][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][442][0]=80'h000000009759c188b4fd;
sos_loop[0].somModel.tcam_mask[6][442][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][443][0]=80'h00000000a08c0f3399b6;
sos_loop[0].somModel.tcam_mask[6][443][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][444][0]=80'h00000000820dea118ef9;
sos_loop[0].somModel.tcam_mask[6][444][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][445][0]=80'h00000000786f4fec3569;
sos_loop[0].somModel.tcam_mask[6][445][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][446][0]=80'h0000000035502a9bf339;
sos_loop[0].somModel.tcam_mask[6][446][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][447][0]=80'h00000000ede032f81911;
sos_loop[0].somModel.tcam_mask[6][447][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][448][0]=80'h00000000005d2da41d57;
sos_loop[0].somModel.tcam_mask[6][448][0]=80'hffffffffff8000000000;
sos_loop[0].somModel.tcam_data[6][449][0]=80'h000000001d551e45233a;
sos_loop[0].somModel.tcam_mask[6][449][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][450][0]=80'h000000001232e7e21619;
sos_loop[0].somModel.tcam_mask[6][450][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][451][0]=80'h000000009656bf8e0b9d;
sos_loop[0].somModel.tcam_mask[6][451][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][452][0]=80'h00000000282df63c9a42;
sos_loop[0].somModel.tcam_mask[6][452][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][453][0]=80'h00000000fb8cfa3efc1a;
sos_loop[0].somModel.tcam_mask[6][453][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][454][0]=80'h00000000e202a5e04142;
sos_loop[0].somModel.tcam_mask[6][454][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][455][0]=80'h00000000ce14bd93ed55;
sos_loop[0].somModel.tcam_mask[6][455][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][456][0]=80'h000000000b29b6b75332;
sos_loop[0].somModel.tcam_mask[6][456][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][457][0]=80'h00000000a560cfe7acfc;
sos_loop[0].somModel.tcam_mask[6][457][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][458][0]=80'h0000000099c7f0448e01;
sos_loop[0].somModel.tcam_mask[6][458][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][459][0]=80'h000000001dc007e9c85a;
sos_loop[0].somModel.tcam_mask[6][459][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][460][0]=80'h00000000d5bbfcebded1;
sos_loop[0].somModel.tcam_mask[6][460][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][461][0]=80'h000000007a59ce859cc7;
sos_loop[0].somModel.tcam_mask[6][461][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][462][0]=80'h000000004ea8c5b70bda;
sos_loop[0].somModel.tcam_mask[6][462][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][463][0]=80'h0000000052f1807fc08a;
sos_loop[0].somModel.tcam_mask[6][463][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][464][0]=80'h00000000206171d9529a;
sos_loop[0].somModel.tcam_mask[6][464][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][465][0]=80'h00000000498a7ea9d6a4;
sos_loop[0].somModel.tcam_mask[6][465][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][466][0]=80'h0000000068b1d8990008;
sos_loop[0].somModel.tcam_mask[6][466][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][467][0]=80'h00000000dfdd7f5c6649;
sos_loop[0].somModel.tcam_mask[6][467][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][468][0]=80'h00000000423c83f43d47;
sos_loop[0].somModel.tcam_mask[6][468][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][469][0]=80'h0000000071daa74440c3;
sos_loop[0].somModel.tcam_mask[6][469][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][470][0]=80'h000000006b7caeb2cb69;
sos_loop[0].somModel.tcam_mask[6][470][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][471][0]=80'h000000009301716b199f;
sos_loop[0].somModel.tcam_mask[6][471][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][472][0]=80'h00000000f30c2c261355;
sos_loop[0].somModel.tcam_mask[6][472][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][473][0]=80'h00000000e1037b5789b6;
sos_loop[0].somModel.tcam_mask[6][473][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][474][0]=80'h000000004ac85c163c30;
sos_loop[0].somModel.tcam_mask[6][474][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][475][0]=80'h00000000bd2e17a3bd71;
sos_loop[0].somModel.tcam_mask[6][475][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][476][0]=80'h000000008cfbaac12a25;
sos_loop[0].somModel.tcam_mask[6][476][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][477][0]=80'h00000000e07f86b355a4;
sos_loop[0].somModel.tcam_mask[6][477][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][478][0]=80'h00000000e24b3b5f435d;
sos_loop[0].somModel.tcam_mask[6][478][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][479][0]=80'h00000000c6100a3221e3;
sos_loop[0].somModel.tcam_mask[6][479][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][480][0]=80'h00000000d601e9e5d6ac;
sos_loop[0].somModel.tcam_mask[6][480][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][481][0]=80'h00000000a2ee82f9007b;
sos_loop[0].somModel.tcam_mask[6][481][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][482][0]=80'h00000000b4baf8944204;
sos_loop[0].somModel.tcam_mask[6][482][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][483][0]=80'h0000000078c5ee1f506d;
sos_loop[0].somModel.tcam_mask[6][483][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][484][0]=80'h0000000094176a64d950;
sos_loop[0].somModel.tcam_mask[6][484][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][485][0]=80'h00000000bdc7edf2bed3;
sos_loop[0].somModel.tcam_mask[6][485][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][486][0]=80'h00000000f6141087125a;
sos_loop[0].somModel.tcam_mask[6][486][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][487][0]=80'h000000004d8a6c4bb175;
sos_loop[0].somModel.tcam_mask[6][487][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][488][0]=80'h00000000d702b7ff755e;
sos_loop[0].somModel.tcam_mask[6][488][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][489][0]=80'h0000000017ad459c4491;
sos_loop[0].somModel.tcam_mask[6][489][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][490][0]=80'h00000000becd69de0af5;
sos_loop[0].somModel.tcam_mask[6][490][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][491][0]=80'h000000006db83a09cb40;
sos_loop[0].somModel.tcam_mask[6][491][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][492][0]=80'h00000000c15a3192c54e;
sos_loop[0].somModel.tcam_mask[6][492][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][493][0]=80'h00000000372729de79a7;
sos_loop[0].somModel.tcam_mask[6][493][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][494][0]=80'h00000000b7d5a573112e;
sos_loop[0].somModel.tcam_mask[6][494][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][495][0]=80'h00000000e7598a8d64ef;
sos_loop[0].somModel.tcam_mask[6][495][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][496][0]=80'h000000004d77a8f186e8;
sos_loop[0].somModel.tcam_mask[6][496][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][497][0]=80'h00000000b3a7e8c62438;
sos_loop[0].somModel.tcam_mask[6][497][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][498][0]=80'h000000005e628e40bad8;
sos_loop[0].somModel.tcam_mask[6][498][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][499][0]=80'h000000002c6ae9566a81;
sos_loop[0].somModel.tcam_mask[6][499][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][500][0]=80'h000000007c8088a4d780;
sos_loop[0].somModel.tcam_mask[6][500][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][501][0]=80'h00000000449da718991b;
sos_loop[0].somModel.tcam_mask[6][501][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][502][0]=80'h00000000eb14915c851e;
sos_loop[0].somModel.tcam_mask[6][502][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][503][0]=80'h000000003527b3d245b5;
sos_loop[0].somModel.tcam_mask[6][503][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][504][0]=80'h0000000085d7cc131a8a;
sos_loop[0].somModel.tcam_mask[6][504][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][505][0]=80'h00000000b448dcc734b3;
sos_loop[0].somModel.tcam_mask[6][505][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][506][0]=80'h000000000463282aaf56;
sos_loop[0].somModel.tcam_mask[6][506][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][507][0]=80'h00000000e6f6fe35b667;
sos_loop[0].somModel.tcam_mask[6][507][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][508][0]=80'h0000000080c258b15826;
sos_loop[0].somModel.tcam_mask[6][508][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][509][0]=80'h00000000faac4f7283f1;
sos_loop[0].somModel.tcam_mask[6][509][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][510][0]=80'h00000000a03cce697a88;
sos_loop[0].somModel.tcam_mask[6][510][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][511][0]=80'h00000000df03c7e186d0;
sos_loop[0].somModel.tcam_mask[6][511][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][512][0]=80'h00000000c301b2ddb491;
sos_loop[0].somModel.tcam_mask[6][512][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][513][0]=80'h0000000005a553a6d946;
sos_loop[0].somModel.tcam_mask[6][513][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][514][0]=80'h00000000ec81a0ecf565;
sos_loop[0].somModel.tcam_mask[6][514][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][515][0]=80'h0000000025b7ba6c7a22;
sos_loop[0].somModel.tcam_mask[6][515][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][516][0]=80'h00000000ff62f77af68e;
sos_loop[0].somModel.tcam_mask[6][516][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][517][0]=80'h0000000090696c0e7c49;
sos_loop[0].somModel.tcam_mask[6][517][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][518][0]=80'h00000000db542752b51b;
sos_loop[0].somModel.tcam_mask[6][518][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][519][0]=80'h000000005c669d7e5719;
sos_loop[0].somModel.tcam_mask[6][519][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][520][0]=80'h0000000007869b90d6d6;
sos_loop[0].somModel.tcam_mask[6][520][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][521][0]=80'h000000006ab3f4028bc4;
sos_loop[0].somModel.tcam_mask[6][521][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][522][0]=80'h00000000faf254c81784;
sos_loop[0].somModel.tcam_mask[6][522][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][523][0]=80'h00000000e91e80ddf2b6;
sos_loop[0].somModel.tcam_mask[6][523][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][524][0]=80'h0000000012ec8002dccf;
sos_loop[0].somModel.tcam_mask[6][524][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][525][0]=80'h000000001fb66119b301;
sos_loop[0].somModel.tcam_mask[6][525][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][526][0]=80'h0000000035cfa56dca6a;
sos_loop[0].somModel.tcam_mask[6][526][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][527][0]=80'h00000000257f17287640;
sos_loop[0].somModel.tcam_mask[6][527][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][528][0]=80'h00000000e24b719e5fd5;
sos_loop[0].somModel.tcam_mask[6][528][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][529][0]=80'h000000001b6de98d63bb;
sos_loop[0].somModel.tcam_mask[6][529][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][530][0]=80'h00000000c7396a1e1d0b;
sos_loop[0].somModel.tcam_mask[6][530][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][531][0]=80'h000000007fb43ae9cd4b;
sos_loop[0].somModel.tcam_mask[6][531][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][532][0]=80'h00000000a389a8825008;
sos_loop[0].somModel.tcam_mask[6][532][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][533][0]=80'h0000000062002cc089d3;
sos_loop[0].somModel.tcam_mask[6][533][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][534][0]=80'h00000000a2fc3e097fd8;
sos_loop[0].somModel.tcam_mask[6][534][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][535][0]=80'h0000000093938f2e7bb6;
sos_loop[0].somModel.tcam_mask[6][535][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][536][0]=80'h000000004c0878c8f3c9;
sos_loop[0].somModel.tcam_mask[6][536][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][537][0]=80'h000000006dad4681d74b;
sos_loop[0].somModel.tcam_mask[6][537][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][538][0]=80'h0000000090d849afd440;
sos_loop[0].somModel.tcam_mask[6][538][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][539][0]=80'h0000000099cea5c192b2;
sos_loop[0].somModel.tcam_mask[6][539][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][540][0]=80'h00000000439a63924ef9;
sos_loop[0].somModel.tcam_mask[6][540][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][541][0]=80'h0000000022efe4c3db4e;
sos_loop[0].somModel.tcam_mask[6][541][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][542][0]=80'h00000000935f8ae1eaca;
sos_loop[0].somModel.tcam_mask[6][542][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][543][0]=80'h00000000980ce89cb3ca;
sos_loop[0].somModel.tcam_mask[6][543][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][544][0]=80'h00000000b2b1d54e6143;
sos_loop[0].somModel.tcam_mask[6][544][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][545][0]=80'h00000000985262ca09c2;
sos_loop[0].somModel.tcam_mask[6][545][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][546][0]=80'h000000001b5370c23148;
sos_loop[0].somModel.tcam_mask[6][546][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][547][0]=80'h00000000fa6e44897737;
sos_loop[0].somModel.tcam_mask[6][547][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][548][0]=80'h00000000edc347b5f551;
sos_loop[0].somModel.tcam_mask[6][548][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][549][0]=80'h00000000bbafbcb86844;
sos_loop[0].somModel.tcam_mask[6][549][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][550][0]=80'h000000007fb9ba95cb59;
sos_loop[0].somModel.tcam_mask[6][550][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][551][0]=80'h00000000be931b35ee21;
sos_loop[0].somModel.tcam_mask[6][551][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][552][0]=80'h0000000039f56d709e34;
sos_loop[0].somModel.tcam_mask[6][552][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][553][0]=80'h000000004e9dfa08200a;
sos_loop[0].somModel.tcam_mask[6][553][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][554][0]=80'h00000000820c31b21a45;
sos_loop[0].somModel.tcam_mask[6][554][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][555][0]=80'h0000000005c7809f7005;
sos_loop[0].somModel.tcam_mask[6][555][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][556][0]=80'h000000003aca0c094cca;
sos_loop[0].somModel.tcam_mask[6][556][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][557][0]=80'h00000000745ae42f60b0;
sos_loop[0].somModel.tcam_mask[6][557][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][558][0]=80'h000000009ab1034e7c6e;
sos_loop[0].somModel.tcam_mask[6][558][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][559][0]=80'h000000008b03e00b02c2;
sos_loop[0].somModel.tcam_mask[6][559][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][560][0]=80'h00000000291393c268aa;
sos_loop[0].somModel.tcam_mask[6][560][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][561][0]=80'h000000004f5dda910b46;
sos_loop[0].somModel.tcam_mask[6][561][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][562][0]=80'h000000000d702572b740;
sos_loop[0].somModel.tcam_mask[6][562][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][563][0]=80'h0000000082eb751a50eb;
sos_loop[0].somModel.tcam_mask[6][563][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][564][0]=80'h0000000069f1bf212be5;
sos_loop[0].somModel.tcam_mask[6][564][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][565][0]=80'h00000000692f8eeae2e9;
sos_loop[0].somModel.tcam_mask[6][565][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][566][0]=80'h0000000019a683169415;
sos_loop[0].somModel.tcam_mask[6][566][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][567][0]=80'h0000000093bac3e6e685;
sos_loop[0].somModel.tcam_mask[6][567][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][568][0]=80'h000000004993bee769ac;
sos_loop[0].somModel.tcam_mask[6][568][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][569][0]=80'h00000000cd7fb4cb6753;
sos_loop[0].somModel.tcam_mask[6][569][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][570][0]=80'h000000000240e7a3c36d;
sos_loop[0].somModel.tcam_mask[6][570][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[6][571][0]=80'h00000000dee7cb29be85;
sos_loop[0].somModel.tcam_mask[6][571][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][572][0]=80'h00000000992597565e42;
sos_loop[0].somModel.tcam_mask[6][572][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][573][0]=80'h000000005cf48819c736;
sos_loop[0].somModel.tcam_mask[6][573][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][574][0]=80'h0000000047abe210da7f;
sos_loop[0].somModel.tcam_mask[6][574][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][575][0]=80'h00000000f93a1757baa0;
sos_loop[0].somModel.tcam_mask[6][575][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][576][0]=80'h000000007c1ceb4afc56;
sos_loop[0].somModel.tcam_mask[6][576][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][577][0]=80'h00000000af7d256d7cc4;
sos_loop[0].somModel.tcam_mask[6][577][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][578][0]=80'h0000000056f4eacb32c7;
sos_loop[0].somModel.tcam_mask[6][578][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][579][0]=80'h00000000b0d1add53e47;
sos_loop[0].somModel.tcam_mask[6][579][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][580][0]=80'h00000000d2755cc4bd17;
sos_loop[0].somModel.tcam_mask[6][580][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][581][0]=80'h00000000a6985589f9f2;
sos_loop[0].somModel.tcam_mask[6][581][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][582][0]=80'h00000000c617a79d7ece;
sos_loop[0].somModel.tcam_mask[6][582][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][583][0]=80'h00000000ce74602fffba;
sos_loop[0].somModel.tcam_mask[6][583][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][584][0]=80'h00000000f924b4b96d61;
sos_loop[0].somModel.tcam_mask[6][584][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][585][0]=80'h000000008c0b6b9901dc;
sos_loop[0].somModel.tcam_mask[6][585][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][586][0]=80'h00000000f68af87708bf;
sos_loop[0].somModel.tcam_mask[6][586][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][587][0]=80'h0000000074fa5f30fe3f;
sos_loop[0].somModel.tcam_mask[6][587][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][588][0]=80'h000000004db8a921b1d2;
sos_loop[0].somModel.tcam_mask[6][588][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][589][0]=80'h0000000018a72f979e24;
sos_loop[0].somModel.tcam_mask[6][589][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][590][0]=80'h00000000595e18260e26;
sos_loop[0].somModel.tcam_mask[6][590][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][591][0]=80'h00000000aad2d483e822;
sos_loop[0].somModel.tcam_mask[6][591][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][592][0]=80'h00000000343913fad305;
sos_loop[0].somModel.tcam_mask[6][592][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][593][0]=80'h00000000b3d2b6c10e97;
sos_loop[0].somModel.tcam_mask[6][593][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][594][0]=80'h000000005b359f4f70b0;
sos_loop[0].somModel.tcam_mask[6][594][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][595][0]=80'h00000000910fdf65238e;
sos_loop[0].somModel.tcam_mask[6][595][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][596][0]=80'h00000000858d2a03d342;
sos_loop[0].somModel.tcam_mask[6][596][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][597][0]=80'h0000000060c0b6079327;
sos_loop[0].somModel.tcam_mask[6][597][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][598][0]=80'h00000000ac7bf03559d7;
sos_loop[0].somModel.tcam_mask[6][598][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][599][0]=80'h000000009ad2390bbe32;
sos_loop[0].somModel.tcam_mask[6][599][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][600][0]=80'h00000000fa4f7ce06718;
sos_loop[0].somModel.tcam_mask[6][600][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][601][0]=80'h00000000d16fe65ec39f;
sos_loop[0].somModel.tcam_mask[6][601][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][602][0]=80'h000000002d99e55053a9;
sos_loop[0].somModel.tcam_mask[6][602][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][603][0]=80'h000000005159029f3697;
sos_loop[0].somModel.tcam_mask[6][603][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][604][0]=80'h00000000b4b0447b5549;
sos_loop[0].somModel.tcam_mask[6][604][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][605][0]=80'h00000000377b752a37b6;
sos_loop[0].somModel.tcam_mask[6][605][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][606][0]=80'h00000000220bb11437f4;
sos_loop[0].somModel.tcam_mask[6][606][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][607][0]=80'h00000000abd69fb1204e;
sos_loop[0].somModel.tcam_mask[6][607][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][608][0]=80'h00000000eb47988d0d8b;
sos_loop[0].somModel.tcam_mask[6][608][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][609][0]=80'h00000000ca9cc767edce;
sos_loop[0].somModel.tcam_mask[6][609][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][610][0]=80'h000000003b6f42cbe0a9;
sos_loop[0].somModel.tcam_mask[6][610][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][611][0]=80'h000000001dd3fa287076;
sos_loop[0].somModel.tcam_mask[6][611][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][612][0]=80'h000000009628912dbff2;
sos_loop[0].somModel.tcam_mask[6][612][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][613][0]=80'h0000000089a7951bea35;
sos_loop[0].somModel.tcam_mask[6][613][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][614][0]=80'h00000000c7b2ff90ab75;
sos_loop[0].somModel.tcam_mask[6][614][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][615][0]=80'h000000007ec37d3f35d1;
sos_loop[0].somModel.tcam_mask[6][615][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][616][0]=80'h00000000486d45350ba4;
sos_loop[0].somModel.tcam_mask[6][616][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][617][0]=80'h00000000f7c78a4aeffd;
sos_loop[0].somModel.tcam_mask[6][617][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][618][0]=80'h00000000ea7f3c4470a0;
sos_loop[0].somModel.tcam_mask[6][618][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][619][0]=80'h0000000095398bca46db;
sos_loop[0].somModel.tcam_mask[6][619][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][620][0]=80'h0000000002a21d269ef9;
sos_loop[0].somModel.tcam_mask[6][620][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[6][621][0]=80'h000000005ff142432afa;
sos_loop[0].somModel.tcam_mask[6][621][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][622][0]=80'h000000008d346fc65e2b;
sos_loop[0].somModel.tcam_mask[6][622][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][623][0]=80'h000000001a6584f50556;
sos_loop[0].somModel.tcam_mask[6][623][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][624][0]=80'h0000000008386da1029f;
sos_loop[0].somModel.tcam_mask[6][624][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][625][0]=80'h00000000db56c981ece6;
sos_loop[0].somModel.tcam_mask[6][625][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][626][0]=80'h00000000cfe8af38f522;
sos_loop[0].somModel.tcam_mask[6][626][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][627][0]=80'h000000008e919d8a745b;
sos_loop[0].somModel.tcam_mask[6][627][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][628][0]=80'h00000000543818958c78;
sos_loop[0].somModel.tcam_mask[6][628][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][629][0]=80'h00000000a8b931f97188;
sos_loop[0].somModel.tcam_mask[6][629][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][630][0]=80'h000000007dee0d849922;
sos_loop[0].somModel.tcam_mask[6][630][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][631][0]=80'h000000001017ca8a2953;
sos_loop[0].somModel.tcam_mask[6][631][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][632][0]=80'h000000007ed9cae24403;
sos_loop[0].somModel.tcam_mask[6][632][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][633][0]=80'h00000000ea187ed4d55a;
sos_loop[0].somModel.tcam_mask[6][633][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][634][0]=80'h000000002e76e28270f1;
sos_loop[0].somModel.tcam_mask[6][634][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][635][0]=80'h00000000f1980343333f;
sos_loop[0].somModel.tcam_mask[6][635][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][636][0]=80'h000000008de1c963c062;
sos_loop[0].somModel.tcam_mask[6][636][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][637][0]=80'h000000003fd86ea44501;
sos_loop[0].somModel.tcam_mask[6][637][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][638][0]=80'h00000000dc791a00bf2c;
sos_loop[0].somModel.tcam_mask[6][638][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][639][0]=80'h0000000076fd772b3105;
sos_loop[0].somModel.tcam_mask[6][639][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][640][0]=80'h000000009137a6d429b2;
sos_loop[0].somModel.tcam_mask[6][640][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][641][0]=80'h0000000049d4cbef7ccc;
sos_loop[0].somModel.tcam_mask[6][641][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][642][0]=80'h000000008051f12b529f;
sos_loop[0].somModel.tcam_mask[6][642][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][643][0]=80'h0000000008d6aa657a5e;
sos_loop[0].somModel.tcam_mask[6][643][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][644][0]=80'h0000000044bafb829ee6;
sos_loop[0].somModel.tcam_mask[6][644][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][645][0]=80'h00000000e55061ccc7b7;
sos_loop[0].somModel.tcam_mask[6][645][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][646][0]=80'h00000000d75970bd3bb0;
sos_loop[0].somModel.tcam_mask[6][646][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][647][0]=80'h000000004811729ba385;
sos_loop[0].somModel.tcam_mask[6][647][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][648][0]=80'h00000000c0501fd955df;
sos_loop[0].somModel.tcam_mask[6][648][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][649][0]=80'h00000000659c29b06d69;
sos_loop[0].somModel.tcam_mask[6][649][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][650][0]=80'h000000006aec373261a3;
sos_loop[0].somModel.tcam_mask[6][650][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][651][0]=80'h00000000c25cd90f5dab;
sos_loop[0].somModel.tcam_mask[6][651][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][652][0]=80'h00000000cee3230bfef6;
sos_loop[0].somModel.tcam_mask[6][652][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][653][0]=80'h000000007bde198a992f;
sos_loop[0].somModel.tcam_mask[6][653][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][654][0]=80'h000000007cd4d9587ccb;
sos_loop[0].somModel.tcam_mask[6][654][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][655][0]=80'h000000005cee7e94dd42;
sos_loop[0].somModel.tcam_mask[6][655][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][656][0]=80'h000000000c7f2c96b613;
sos_loop[0].somModel.tcam_mask[6][656][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][657][0]=80'h00000000f2de9d0bdde4;
sos_loop[0].somModel.tcam_mask[6][657][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][658][0]=80'h00000000b80342294761;
sos_loop[0].somModel.tcam_mask[6][658][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][659][0]=80'h00000000ef05f9051dde;
sos_loop[0].somModel.tcam_mask[6][659][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][660][0]=80'h00000000089d9864b0f7;
sos_loop[0].somModel.tcam_mask[6][660][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[6][661][0]=80'h00000000f84ebc6b5933;
sos_loop[0].somModel.tcam_mask[6][661][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][662][0]=80'h0000000099c7ebd6ef11;
sos_loop[0].somModel.tcam_mask[6][662][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][663][0]=80'h00000000a5cfc726453c;
sos_loop[0].somModel.tcam_mask[6][663][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][664][0]=80'h000000008e33ccc43905;
sos_loop[0].somModel.tcam_mask[6][664][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][665][0]=80'h0000000061dbc393f8b8;
sos_loop[0].somModel.tcam_mask[6][665][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][666][0]=80'h00000000b5776eb8e40c;
sos_loop[0].somModel.tcam_mask[6][666][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][667][0]=80'h00000000c56f02fbb8af;
sos_loop[0].somModel.tcam_mask[6][667][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][668][0]=80'h00000000f06ac89a6e2e;
sos_loop[0].somModel.tcam_mask[6][668][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][669][0]=80'h000000004d46ea5704c7;
sos_loop[0].somModel.tcam_mask[6][669][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][670][0]=80'h00000000018a0d2ab536;
sos_loop[0].somModel.tcam_mask[6][670][0]=80'hfffffffffe0000000000;
sos_loop[0].somModel.tcam_data[6][671][0]=80'h00000000de24ea9c8559;
sos_loop[0].somModel.tcam_mask[6][671][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][672][0]=80'h00000000117c2dcb8a3f;
sos_loop[0].somModel.tcam_mask[6][672][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][673][0]=80'h00000000042c5800a198;
sos_loop[0].somModel.tcam_mask[6][673][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][674][0]=80'h00000000c866641162c8;
sos_loop[0].somModel.tcam_mask[6][674][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][675][0]=80'h00000000c59ce2a178ef;
sos_loop[0].somModel.tcam_mask[6][675][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][676][0]=80'h0000000091b9a88b2186;
sos_loop[0].somModel.tcam_mask[6][676][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][677][0]=80'h00000000baaaa92f9330;
sos_loop[0].somModel.tcam_mask[6][677][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][678][0]=80'h00000000899bc4d45fed;
sos_loop[0].somModel.tcam_mask[6][678][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][679][0]=80'h0000000031aba86c07cd;
sos_loop[0].somModel.tcam_mask[6][679][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][680][0]=80'h00000000c4984e56b9a3;
sos_loop[0].somModel.tcam_mask[6][680][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][681][0]=80'h000000001b2cb5378bd2;
sos_loop[0].somModel.tcam_mask[6][681][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[6][682][0]=80'h00000000ff120ca68f9a;
sos_loop[0].somModel.tcam_mask[6][682][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][683][0]=80'h00000000a835dfd4a64e;
sos_loop[0].somModel.tcam_mask[6][683][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][684][0]=80'h00000000cc35683c57dc;
sos_loop[0].somModel.tcam_mask[6][684][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][685][0]=80'h00000000a5c1099a0ccc;
sos_loop[0].somModel.tcam_mask[6][685][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][686][0]=80'h00000000efd95c4e5fe9;
sos_loop[0].somModel.tcam_mask[6][686][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][687][0]=80'h000000007c76d25796aa;
sos_loop[0].somModel.tcam_mask[6][687][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][688][0]=80'h0000000007b60730923d;
sos_loop[0].somModel.tcam_mask[6][688][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][689][0]=80'h0000000007373b8b8f3c;
sos_loop[0].somModel.tcam_mask[6][689][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[6][690][0]=80'h0000000037e56c799b77;
sos_loop[0].somModel.tcam_mask[6][690][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[6][691][0]=80'h0000000064aeec7ab84c;
sos_loop[0].somModel.tcam_mask[6][691][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][692][0]=80'h00000000dc1814387312;
sos_loop[0].somModel.tcam_mask[6][692][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][693][0]=80'h00000000dd2835b8c4f9;
sos_loop[0].somModel.tcam_mask[6][693][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][694][0]=80'h000000005af2eb552cca;
sos_loop[0].somModel.tcam_mask[6][694][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][695][0]=80'h00000000446b9299fa74;
sos_loop[0].somModel.tcam_mask[6][695][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][696][0]=80'h0000000086928cf64fc6;
sos_loop[0].somModel.tcam_mask[6][696][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][697][0]=80'h00000000c4fdc019c61f;
sos_loop[0].somModel.tcam_mask[6][697][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][698][0]=80'h00000000882f97bb161f;
sos_loop[0].somModel.tcam_mask[6][698][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[6][699][0]=80'h000000004ed606f4518d;
sos_loop[0].somModel.tcam_mask[6][699][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[6][700][0]=80'h00000000bd46a3aa3c15;
sos_loop[0].somModel.tcam_mask[6][700][0]=80'hffffffff000000000000;
sos_loop[0].somModel.sram_dat[6][0][0]=96'hdeadbf;
sos_loop[0].somModel.sram_ptr[6][0]=939;
sos_loop[0].somModel.sram_dat[6][1][0]=96'hc153;
sos_loop[0].somModel.sram_ptr[6][1]=3;
sos_loop[0].somModel.sram_dat[6][2][0]=96'hdf3d;
sos_loop[0].somModel.sram_ptr[6][2]=3;
sos_loop[0].somModel.sram_dat[6][3][0]=96'h3f56;
sos_loop[0].somModel.sram_ptr[6][3]=3;
sos_loop[0].somModel.sram_dat[6][4][0]=96'hb758;
sos_loop[0].somModel.sram_ptr[6][4]=3;
sos_loop[0].somModel.sram_dat[6][5][0]=96'h972b;
sos_loop[0].somModel.sram_ptr[6][5]=3;
sos_loop[0].somModel.sram_dat[6][6][0]=96'h624e;
sos_loop[0].somModel.sram_ptr[6][6]=3;
sos_loop[0].somModel.sram_dat[6][7][0]=96'hd51d;
sos_loop[0].somModel.sram_ptr[6][7]=3;
sos_loop[0].somModel.sram_dat[6][8][0]=96'hb905;
sos_loop[0].somModel.sram_ptr[6][8]=3;
sos_loop[0].somModel.sram_dat[6][9][0]=96'ha8a9;
sos_loop[0].somModel.sram_ptr[6][9]=3;
sos_loop[0].somModel.sram_dat[6][10][0]=96'ha7c9;
sos_loop[0].somModel.sram_ptr[6][10]=3;
sos_loop[0].somModel.sram_dat[6][11][0]=96'h37f8;
sos_loop[0].somModel.sram_ptr[6][11]=3;
sos_loop[0].somModel.sram_dat[6][12][0]=96'hee8c;
sos_loop[0].somModel.sram_ptr[6][12]=3;
sos_loop[0].somModel.sram_dat[6][13][0]=96'h95f5;
sos_loop[0].somModel.sram_ptr[6][13]=3;
sos_loop[0].somModel.sram_dat[6][14][0]=96'hbe40;
sos_loop[0].somModel.sram_ptr[6][14]=3;
sos_loop[0].somModel.sram_dat[6][15][0]=96'ha2c3;
sos_loop[0].somModel.sram_ptr[6][15]=3;
sos_loop[0].somModel.sram_dat[6][16][0]=96'h3275;
sos_loop[0].somModel.sram_ptr[6][16]=3;
sos_loop[0].somModel.sram_dat[6][17][0]=96'hf5ff;
sos_loop[0].somModel.sram_ptr[6][17]=3;
sos_loop[0].somModel.sram_dat[6][18][0]=96'h84c6;
sos_loop[0].somModel.sram_ptr[6][18]=3;
sos_loop[0].somModel.sram_dat[6][19][0]=96'ha54c;
sos_loop[0].somModel.sram_ptr[6][19]=3;
sos_loop[0].somModel.sram_dat[6][20][0]=96'hc4f3;
sos_loop[0].somModel.sram_ptr[6][20]=3;
sos_loop[0].somModel.sram_dat[6][21][0]=96'h4a8d;
sos_loop[0].somModel.sram_ptr[6][21]=3;
sos_loop[0].somModel.sram_dat[6][22][0]=96'hfe35;
sos_loop[0].somModel.sram_ptr[6][22]=3;
sos_loop[0].somModel.sram_dat[6][23][0]=96'hdff6;
sos_loop[0].somModel.sram_ptr[6][23]=3;
sos_loop[0].somModel.sram_dat[6][24][0]=96'h1765;
sos_loop[0].somModel.sram_ptr[6][24]=3;
sos_loop[0].somModel.sram_dat[6][25][0]=96'hb292;
sos_loop[0].somModel.sram_ptr[6][25]=3;
sos_loop[0].somModel.sram_dat[6][26][0]=96'h4d71;
sos_loop[0].somModel.sram_ptr[6][26]=3;
sos_loop[0].somModel.sram_dat[6][27][0]=96'h4d83;
sos_loop[0].somModel.sram_ptr[6][27]=3;
sos_loop[0].somModel.sram_dat[6][28][0]=96'h6c69;
sos_loop[0].somModel.sram_ptr[6][28]=3;
sos_loop[0].somModel.sram_dat[6][29][0]=96'h1c6b;
sos_loop[0].somModel.sram_ptr[6][29]=3;
sos_loop[0].somModel.sram_dat[6][30][0]=96'ha4bb;
sos_loop[0].somModel.sram_ptr[6][30]=3;
sos_loop[0].somModel.sram_dat[6][31][0]=96'h9c42;
sos_loop[0].somModel.sram_ptr[6][31]=3;
sos_loop[0].somModel.sram_dat[6][32][0]=96'hf399;
sos_loop[0].somModel.sram_ptr[6][32]=3;
sos_loop[0].somModel.sram_dat[6][33][0]=96'he276;
sos_loop[0].somModel.sram_ptr[6][33]=3;
sos_loop[0].somModel.sram_dat[6][34][0]=96'h782c;
sos_loop[0].somModel.sram_ptr[6][34]=3;
sos_loop[0].somModel.sram_dat[6][35][0]=96'h556;
sos_loop[0].somModel.sram_ptr[6][35]=3;
sos_loop[0].somModel.sram_dat[6][36][0]=96'h3d19;
sos_loop[0].somModel.sram_ptr[6][36]=3;
sos_loop[0].somModel.sram_dat[6][37][0]=96'h61df;
sos_loop[0].somModel.sram_ptr[6][37]=3;
sos_loop[0].somModel.sram_dat[6][38][0]=96'h25c0;
sos_loop[0].somModel.sram_ptr[6][38]=3;
sos_loop[0].somModel.sram_dat[6][39][0]=96'h4c4b;
sos_loop[0].somModel.sram_ptr[6][39]=3;
sos_loop[0].somModel.sram_dat[6][40][0]=96'h962;
sos_loop[0].somModel.sram_ptr[6][40]=3;
sos_loop[0].somModel.sram_dat[6][41][0]=96'ha4e4;
sos_loop[0].somModel.sram_ptr[6][41]=3;
sos_loop[0].somModel.sram_dat[6][42][0]=96'h3376;
sos_loop[0].somModel.sram_ptr[6][42]=3;
sos_loop[0].somModel.sram_dat[6][43][0]=96'hbfd6;
sos_loop[0].somModel.sram_ptr[6][43]=3;
sos_loop[0].somModel.sram_dat[6][44][0]=96'h2121;
sos_loop[0].somModel.sram_ptr[6][44]=3;
sos_loop[0].somModel.sram_dat[6][45][0]=96'h393a;
sos_loop[0].somModel.sram_ptr[6][45]=3;
sos_loop[0].somModel.sram_dat[6][46][0]=96'hc59c;
sos_loop[0].somModel.sram_ptr[6][46]=3;
sos_loop[0].somModel.sram_dat[6][47][0]=96'hbab5;
sos_loop[0].somModel.sram_ptr[6][47]=3;
sos_loop[0].somModel.sram_dat[6][48][0]=96'h4d89;
sos_loop[0].somModel.sram_ptr[6][48]=3;
sos_loop[0].somModel.sram_dat[6][49][0]=96'h78ec;
sos_loop[0].somModel.sram_ptr[6][49]=3;
sos_loop[0].somModel.sram_dat[6][50][0]=96'h9051;
sos_loop[0].somModel.sram_ptr[6][50]=3;
sos_loop[0].somModel.sram_dat[6][51][0]=96'h1fb5;
sos_loop[0].somModel.sram_ptr[6][51]=3;
sos_loop[0].somModel.sram_dat[6][52][0]=96'h84c3;
sos_loop[0].somModel.sram_ptr[6][52]=3;
sos_loop[0].somModel.sram_dat[6][53][0]=96'h532f;
sos_loop[0].somModel.sram_ptr[6][53]=3;
sos_loop[0].somModel.sram_dat[6][54][0]=96'hfcec;
sos_loop[0].somModel.sram_ptr[6][54]=3;
sos_loop[0].somModel.sram_dat[6][55][0]=96'h460e;
sos_loop[0].somModel.sram_ptr[6][55]=3;
sos_loop[0].somModel.sram_dat[6][56][0]=96'h12a9;
sos_loop[0].somModel.sram_ptr[6][56]=3;
sos_loop[0].somModel.sram_dat[6][57][0]=96'h2f22;
sos_loop[0].somModel.sram_ptr[6][57]=3;
sos_loop[0].somModel.sram_dat[6][58][0]=96'h297d;
sos_loop[0].somModel.sram_ptr[6][58]=3;
sos_loop[0].somModel.sram_dat[6][59][0]=96'h2f95;
sos_loop[0].somModel.sram_ptr[6][59]=3;
sos_loop[0].somModel.sram_dat[6][60][0]=96'h3952;
sos_loop[0].somModel.sram_ptr[6][60]=3;
sos_loop[0].somModel.sram_dat[6][61][0]=96'h59e5;
sos_loop[0].somModel.sram_ptr[6][61]=3;
sos_loop[0].somModel.sram_dat[6][62][0]=96'h4201;
sos_loop[0].somModel.sram_ptr[6][62]=3;
sos_loop[0].somModel.sram_dat[6][63][0]=96'habfb;
sos_loop[0].somModel.sram_ptr[6][63]=3;
sos_loop[0].somModel.sram_dat[6][64][0]=96'h890f;
sos_loop[0].somModel.sram_ptr[6][64]=3;
sos_loop[0].somModel.sram_dat[6][65][0]=96'hfc14;
sos_loop[0].somModel.sram_ptr[6][65]=3;
sos_loop[0].somModel.sram_dat[6][66][0]=96'h561d;
sos_loop[0].somModel.sram_ptr[6][66]=3;
sos_loop[0].somModel.sram_dat[6][67][0]=96'h9b06;
sos_loop[0].somModel.sram_ptr[6][67]=3;
sos_loop[0].somModel.sram_dat[6][68][0]=96'hc82;
sos_loop[0].somModel.sram_ptr[6][68]=3;
sos_loop[0].somModel.sram_dat[6][69][0]=96'h7392;
sos_loop[0].somModel.sram_ptr[6][69]=3;
sos_loop[0].somModel.sram_dat[6][70][0]=96'h69f8;
sos_loop[0].somModel.sram_ptr[6][70]=3;
sos_loop[0].somModel.sram_dat[6][71][0]=96'hab52;
sos_loop[0].somModel.sram_ptr[6][71]=3;
sos_loop[0].somModel.sram_dat[6][72][0]=96'h46a7;
sos_loop[0].somModel.sram_ptr[6][72]=3;
sos_loop[0].somModel.sram_dat[6][73][0]=96'h88bd;
sos_loop[0].somModel.sram_ptr[6][73]=3;
sos_loop[0].somModel.sram_dat[6][74][0]=96'hb6c5;
sos_loop[0].somModel.sram_ptr[6][74]=3;
sos_loop[0].somModel.sram_dat[6][75][0]=96'hf611;
sos_loop[0].somModel.sram_ptr[6][75]=3;
sos_loop[0].somModel.sram_dat[6][76][0]=96'h1778;
sos_loop[0].somModel.sram_ptr[6][76]=3;
sos_loop[0].somModel.sram_dat[6][77][0]=96'h9317;
sos_loop[0].somModel.sram_ptr[6][77]=3;
sos_loop[0].somModel.sram_dat[6][78][0]=96'hb32f;
sos_loop[0].somModel.sram_ptr[6][78]=3;
sos_loop[0].somModel.sram_dat[6][79][0]=96'hf584;
sos_loop[0].somModel.sram_ptr[6][79]=3;
sos_loop[0].somModel.sram_dat[6][80][0]=96'h1183;
sos_loop[0].somModel.sram_ptr[6][80]=3;
sos_loop[0].somModel.sram_dat[6][81][0]=96'he56f;
sos_loop[0].somModel.sram_ptr[6][81]=3;
sos_loop[0].somModel.sram_dat[6][82][0]=96'h73f8;
sos_loop[0].somModel.sram_ptr[6][82]=3;
sos_loop[0].somModel.sram_dat[6][83][0]=96'he077;
sos_loop[0].somModel.sram_ptr[6][83]=3;
sos_loop[0].somModel.sram_dat[6][84][0]=96'h9ca6;
sos_loop[0].somModel.sram_ptr[6][84]=3;
sos_loop[0].somModel.sram_dat[6][85][0]=96'h9acc;
sos_loop[0].somModel.sram_ptr[6][85]=3;
sos_loop[0].somModel.sram_dat[6][86][0]=96'h165c;
sos_loop[0].somModel.sram_ptr[6][86]=3;
sos_loop[0].somModel.sram_dat[6][87][0]=96'h956e;
sos_loop[0].somModel.sram_ptr[6][87]=3;
sos_loop[0].somModel.sram_dat[6][88][0]=96'ha541;
sos_loop[0].somModel.sram_ptr[6][88]=3;
sos_loop[0].somModel.sram_dat[6][89][0]=96'hb89e;
sos_loop[0].somModel.sram_ptr[6][89]=3;
sos_loop[0].somModel.sram_dat[6][90][0]=96'h3001;
sos_loop[0].somModel.sram_ptr[6][90]=3;
sos_loop[0].somModel.sram_dat[6][91][0]=96'h23b7;
sos_loop[0].somModel.sram_ptr[6][91]=3;
sos_loop[0].somModel.sram_dat[6][92][0]=96'ha9b2;
sos_loop[0].somModel.sram_ptr[6][92]=3;
sos_loop[0].somModel.sram_dat[6][93][0]=96'hf128;
sos_loop[0].somModel.sram_ptr[6][93]=3;
sos_loop[0].somModel.sram_dat[6][94][0]=96'hb305;
sos_loop[0].somModel.sram_ptr[6][94]=3;
sos_loop[0].somModel.sram_dat[6][95][0]=96'h32;
sos_loop[0].somModel.sram_ptr[6][95]=3;
sos_loop[0].somModel.sram_dat[6][96][0]=96'h1876;
sos_loop[0].somModel.sram_ptr[6][96]=3;
sos_loop[0].somModel.sram_dat[6][97][0]=96'hf881;
sos_loop[0].somModel.sram_ptr[6][97]=3;
sos_loop[0].somModel.sram_dat[6][98][0]=96'hdbfb;
sos_loop[0].somModel.sram_ptr[6][98]=3;
sos_loop[0].somModel.sram_dat[6][99][0]=96'haa91;
sos_loop[0].somModel.sram_ptr[6][99]=3;
sos_loop[0].somModel.sram_dat[6][100][0]=96'h4b52;
sos_loop[0].somModel.sram_ptr[6][100]=3;
sos_loop[0].somModel.sram_dat[6][101][0]=96'hb267;
sos_loop[0].somModel.sram_ptr[6][101]=3;
sos_loop[0].somModel.sram_dat[6][102][0]=96'h7b38;
sos_loop[0].somModel.sram_ptr[6][102]=3;
sos_loop[0].somModel.sram_dat[6][103][0]=96'h3af9;
sos_loop[0].somModel.sram_ptr[6][103]=3;
sos_loop[0].somModel.sram_dat[6][104][0]=96'h1df7;
sos_loop[0].somModel.sram_ptr[6][104]=3;
sos_loop[0].somModel.sram_dat[6][105][0]=96'hf165;
sos_loop[0].somModel.sram_ptr[6][105]=3;
sos_loop[0].somModel.sram_dat[6][106][0]=96'h202f;
sos_loop[0].somModel.sram_ptr[6][106]=3;
sos_loop[0].somModel.sram_dat[6][107][0]=96'h40c4;
sos_loop[0].somModel.sram_ptr[6][107]=3;
sos_loop[0].somModel.sram_dat[6][108][0]=96'h1275;
sos_loop[0].somModel.sram_ptr[6][108]=3;
sos_loop[0].somModel.sram_dat[6][109][0]=96'h67fe;
sos_loop[0].somModel.sram_ptr[6][109]=3;
sos_loop[0].somModel.sram_dat[6][110][0]=96'h23a4;
sos_loop[0].somModel.sram_ptr[6][110]=3;
sos_loop[0].somModel.sram_dat[6][111][0]=96'h311d;
sos_loop[0].somModel.sram_ptr[6][111]=3;
sos_loop[0].somModel.sram_dat[6][112][0]=96'h995f;
sos_loop[0].somModel.sram_ptr[6][112]=3;
sos_loop[0].somModel.sram_dat[6][113][0]=96'h6a35;
sos_loop[0].somModel.sram_ptr[6][113]=3;
sos_loop[0].somModel.sram_dat[6][114][0]=96'hc8;
sos_loop[0].somModel.sram_ptr[6][114]=3;
sos_loop[0].somModel.sram_dat[6][115][0]=96'h3087;
sos_loop[0].somModel.sram_ptr[6][115]=3;
sos_loop[0].somModel.sram_dat[6][116][0]=96'hf1b6;
sos_loop[0].somModel.sram_ptr[6][116]=3;
sos_loop[0].somModel.sram_dat[6][117][0]=96'h7805;
sos_loop[0].somModel.sram_ptr[6][117]=3;
sos_loop[0].somModel.sram_dat[6][118][0]=96'ha535;
sos_loop[0].somModel.sram_ptr[6][118]=3;
sos_loop[0].somModel.sram_dat[6][119][0]=96'hffca;
sos_loop[0].somModel.sram_ptr[6][119]=3;
sos_loop[0].somModel.sram_dat[6][120][0]=96'hfa15;
sos_loop[0].somModel.sram_ptr[6][120]=3;
sos_loop[0].somModel.sram_dat[6][121][0]=96'hde2d;
sos_loop[0].somModel.sram_ptr[6][121]=3;
sos_loop[0].somModel.sram_dat[6][122][0]=96'h2fcb;
sos_loop[0].somModel.sram_ptr[6][122]=3;
sos_loop[0].somModel.sram_dat[6][123][0]=96'h432c;
sos_loop[0].somModel.sram_ptr[6][123]=3;
sos_loop[0].somModel.sram_dat[6][124][0]=96'hf151;
sos_loop[0].somModel.sram_ptr[6][124]=3;
sos_loop[0].somModel.sram_dat[6][125][0]=96'hdd1e;
sos_loop[0].somModel.sram_ptr[6][125]=3;
sos_loop[0].somModel.sram_dat[6][126][0]=96'ha8c6;
sos_loop[0].somModel.sram_ptr[6][126]=3;
sos_loop[0].somModel.sram_dat[6][127][0]=96'h8146;
sos_loop[0].somModel.sram_ptr[6][127]=3;
sos_loop[0].somModel.sram_dat[6][128][0]=96'h86b9;
sos_loop[0].somModel.sram_ptr[6][128]=3;
sos_loop[0].somModel.sram_dat[6][129][0]=96'h6bda;
sos_loop[0].somModel.sram_ptr[6][129]=3;
sos_loop[0].somModel.sram_dat[6][130][0]=96'h35d5;
sos_loop[0].somModel.sram_ptr[6][130]=3;
sos_loop[0].somModel.sram_dat[6][131][0]=96'h7354;
sos_loop[0].somModel.sram_ptr[6][131]=3;
sos_loop[0].somModel.sram_dat[6][132][0]=96'he59b;
sos_loop[0].somModel.sram_ptr[6][132]=3;
sos_loop[0].somModel.sram_dat[6][133][0]=96'h4237;
sos_loop[0].somModel.sram_ptr[6][133]=3;
sos_loop[0].somModel.sram_dat[6][134][0]=96'h4b8c;
sos_loop[0].somModel.sram_ptr[6][134]=3;
sos_loop[0].somModel.sram_dat[6][135][0]=96'h1a7a;
sos_loop[0].somModel.sram_ptr[6][135]=3;
sos_loop[0].somModel.sram_dat[6][136][0]=96'h181b;
sos_loop[0].somModel.sram_ptr[6][136]=3;
sos_loop[0].somModel.sram_dat[6][137][0]=96'h610a;
sos_loop[0].somModel.sram_ptr[6][137]=3;
sos_loop[0].somModel.sram_dat[6][138][0]=96'h6087;
sos_loop[0].somModel.sram_ptr[6][138]=3;
sos_loop[0].somModel.sram_dat[6][139][0]=96'h5869;
sos_loop[0].somModel.sram_ptr[6][139]=3;
sos_loop[0].somModel.sram_dat[6][140][0]=96'h6af7;
sos_loop[0].somModel.sram_ptr[6][140]=3;
sos_loop[0].somModel.sram_dat[6][141][0]=96'h9b7f;
sos_loop[0].somModel.sram_ptr[6][141]=3;
sos_loop[0].somModel.sram_dat[6][142][0]=96'hc12a;
sos_loop[0].somModel.sram_ptr[6][142]=3;
sos_loop[0].somModel.sram_dat[6][143][0]=96'h7112;
sos_loop[0].somModel.sram_ptr[6][143]=3;
sos_loop[0].somModel.sram_dat[6][144][0]=96'hff31;
sos_loop[0].somModel.sram_ptr[6][144]=3;
sos_loop[0].somModel.sram_dat[6][145][0]=96'hb651;
sos_loop[0].somModel.sram_ptr[6][145]=3;
sos_loop[0].somModel.sram_dat[6][146][0]=96'h4243;
sos_loop[0].somModel.sram_ptr[6][146]=3;
sos_loop[0].somModel.sram_dat[6][147][0]=96'hb299;
sos_loop[0].somModel.sram_ptr[6][147]=3;
sos_loop[0].somModel.sram_dat[6][148][0]=96'h7605;
sos_loop[0].somModel.sram_ptr[6][148]=3;
sos_loop[0].somModel.sram_dat[6][149][0]=96'he4a2;
sos_loop[0].somModel.sram_ptr[6][149]=3;
sos_loop[0].somModel.sram_dat[6][150][0]=96'he751;
sos_loop[0].somModel.sram_ptr[6][150]=3;
sos_loop[0].somModel.sram_dat[6][151][0]=96'hedf2;
sos_loop[0].somModel.sram_ptr[6][151]=3;
sos_loop[0].somModel.sram_dat[6][152][0]=96'h3cfc;
sos_loop[0].somModel.sram_ptr[6][152]=3;
sos_loop[0].somModel.sram_dat[6][153][0]=96'hc7ba;
sos_loop[0].somModel.sram_ptr[6][153]=3;
sos_loop[0].somModel.sram_dat[6][154][0]=96'hc156;
sos_loop[0].somModel.sram_ptr[6][154]=3;
sos_loop[0].somModel.sram_dat[6][155][0]=96'h81aa;
sos_loop[0].somModel.sram_ptr[6][155]=3;
sos_loop[0].somModel.sram_dat[6][156][0]=96'he58f;
sos_loop[0].somModel.sram_ptr[6][156]=3;
sos_loop[0].somModel.sram_dat[6][157][0]=96'h8635;
sos_loop[0].somModel.sram_ptr[6][157]=3;
sos_loop[0].somModel.sram_dat[6][158][0]=96'haf80;
sos_loop[0].somModel.sram_ptr[6][158]=3;
sos_loop[0].somModel.sram_dat[6][159][0]=96'hbad8;
sos_loop[0].somModel.sram_ptr[6][159]=3;
sos_loop[0].somModel.sram_dat[6][160][0]=96'hbcfb;
sos_loop[0].somModel.sram_ptr[6][160]=3;
sos_loop[0].somModel.sram_dat[6][161][0]=96'h4b9c;
sos_loop[0].somModel.sram_ptr[6][161]=3;
sos_loop[0].somModel.sram_dat[6][162][0]=96'h72e2;
sos_loop[0].somModel.sram_ptr[6][162]=3;
sos_loop[0].somModel.sram_dat[6][163][0]=96'hc60d;
sos_loop[0].somModel.sram_ptr[6][163]=3;
sos_loop[0].somModel.sram_dat[6][164][0]=96'ha224;
sos_loop[0].somModel.sram_ptr[6][164]=3;
sos_loop[0].somModel.sram_dat[6][165][0]=96'h52f;
sos_loop[0].somModel.sram_ptr[6][165]=3;
sos_loop[0].somModel.sram_dat[6][166][0]=96'h1ede;
sos_loop[0].somModel.sram_ptr[6][166]=3;
sos_loop[0].somModel.sram_dat[6][167][0]=96'h41a4;
sos_loop[0].somModel.sram_ptr[6][167]=3;
sos_loop[0].somModel.sram_dat[6][168][0]=96'h615;
sos_loop[0].somModel.sram_ptr[6][168]=3;
sos_loop[0].somModel.sram_dat[6][169][0]=96'h31b1;
sos_loop[0].somModel.sram_ptr[6][169]=3;
sos_loop[0].somModel.sram_dat[6][170][0]=96'hf78f;
sos_loop[0].somModel.sram_ptr[6][170]=3;
sos_loop[0].somModel.sram_dat[6][171][0]=96'hc802;
sos_loop[0].somModel.sram_ptr[6][171]=3;
sos_loop[0].somModel.sram_dat[6][172][0]=96'h829a;
sos_loop[0].somModel.sram_ptr[6][172]=3;
sos_loop[0].somModel.sram_dat[6][173][0]=96'h3866;
sos_loop[0].somModel.sram_ptr[6][173]=3;
sos_loop[0].somModel.sram_dat[6][174][0]=96'he962;
sos_loop[0].somModel.sram_ptr[6][174]=3;
sos_loop[0].somModel.sram_dat[6][175][0]=96'h12f;
sos_loop[0].somModel.sram_ptr[6][175]=3;
sos_loop[0].somModel.sram_dat[6][176][0]=96'h90b9;
sos_loop[0].somModel.sram_ptr[6][176]=3;
sos_loop[0].somModel.sram_dat[6][177][0]=96'ha9bc;
sos_loop[0].somModel.sram_ptr[6][177]=3;
sos_loop[0].somModel.sram_dat[6][178][0]=96'h8f6d;
sos_loop[0].somModel.sram_ptr[6][178]=3;
sos_loop[0].somModel.sram_dat[6][179][0]=96'h173a;
sos_loop[0].somModel.sram_ptr[6][179]=3;
sos_loop[0].somModel.sram_dat[6][180][0]=96'h204c;
sos_loop[0].somModel.sram_ptr[6][180]=3;
sos_loop[0].somModel.sram_dat[6][181][0]=96'hf907;
sos_loop[0].somModel.sram_ptr[6][181]=3;
sos_loop[0].somModel.sram_dat[6][182][0]=96'hfc36;
sos_loop[0].somModel.sram_ptr[6][182]=3;
sos_loop[0].somModel.sram_dat[6][183][0]=96'hd4c8;
sos_loop[0].somModel.sram_ptr[6][183]=3;
sos_loop[0].somModel.sram_dat[6][184][0]=96'hcff9;
sos_loop[0].somModel.sram_ptr[6][184]=3;
sos_loop[0].somModel.sram_dat[6][185][0]=96'h167e;
sos_loop[0].somModel.sram_ptr[6][185]=3;
sos_loop[0].somModel.sram_dat[6][186][0]=96'hd549;
sos_loop[0].somModel.sram_ptr[6][186]=3;
sos_loop[0].somModel.sram_dat[6][187][0]=96'hef1;
sos_loop[0].somModel.sram_ptr[6][187]=3;
sos_loop[0].somModel.sram_dat[6][188][0]=96'h197;
sos_loop[0].somModel.sram_ptr[6][188]=3;
sos_loop[0].somModel.sram_dat[6][189][0]=96'hd74c;
sos_loop[0].somModel.sram_ptr[6][189]=3;
sos_loop[0].somModel.sram_dat[6][190][0]=96'haa47;
sos_loop[0].somModel.sram_ptr[6][190]=3;
sos_loop[0].somModel.sram_dat[6][191][0]=96'h457b;
sos_loop[0].somModel.sram_ptr[6][191]=3;
sos_loop[0].somModel.sram_dat[6][192][0]=96'he8d2;
sos_loop[0].somModel.sram_ptr[6][192]=3;
sos_loop[0].somModel.sram_dat[6][193][0]=96'h43db;
sos_loop[0].somModel.sram_ptr[6][193]=3;
sos_loop[0].somModel.sram_dat[6][194][0]=96'hb4cd;
sos_loop[0].somModel.sram_ptr[6][194]=3;
sos_loop[0].somModel.sram_dat[6][195][0]=96'h3320;
sos_loop[0].somModel.sram_ptr[6][195]=3;
sos_loop[0].somModel.sram_dat[6][196][0]=96'hf172;
sos_loop[0].somModel.sram_ptr[6][196]=3;
sos_loop[0].somModel.sram_dat[6][197][0]=96'hab6c;
sos_loop[0].somModel.sram_ptr[6][197]=3;
sos_loop[0].somModel.sram_dat[6][198][0]=96'h10d1;
sos_loop[0].somModel.sram_ptr[6][198]=3;
sos_loop[0].somModel.sram_dat[6][199][0]=96'hc1de;
sos_loop[0].somModel.sram_ptr[6][199]=3;
sos_loop[0].somModel.sram_dat[6][200][0]=96'h4a5;
sos_loop[0].somModel.sram_ptr[6][200]=3;
sos_loop[0].somModel.sram_dat[6][201][0]=96'h4677;
sos_loop[0].somModel.sram_ptr[6][201]=3;
sos_loop[0].somModel.sram_dat[6][202][0]=96'h1955;
sos_loop[0].somModel.sram_ptr[6][202]=3;
sos_loop[0].somModel.sram_dat[6][203][0]=96'h2287;
sos_loop[0].somModel.sram_ptr[6][203]=3;
sos_loop[0].somModel.sram_dat[6][204][0]=96'h7fbc;
sos_loop[0].somModel.sram_ptr[6][204]=3;
sos_loop[0].somModel.sram_dat[6][205][0]=96'h5226;
sos_loop[0].somModel.sram_ptr[6][205]=3;
sos_loop[0].somModel.sram_dat[6][206][0]=96'he45e;
sos_loop[0].somModel.sram_ptr[6][206]=3;
sos_loop[0].somModel.sram_dat[6][207][0]=96'hc5d6;
sos_loop[0].somModel.sram_ptr[6][207]=3;
sos_loop[0].somModel.sram_dat[6][208][0]=96'h592e;
sos_loop[0].somModel.sram_ptr[6][208]=3;
sos_loop[0].somModel.sram_dat[6][209][0]=96'he0dd;
sos_loop[0].somModel.sram_ptr[6][209]=3;
sos_loop[0].somModel.sram_dat[6][210][0]=96'h5cd3;
sos_loop[0].somModel.sram_ptr[6][210]=3;
sos_loop[0].somModel.sram_dat[6][211][0]=96'h4976;
sos_loop[0].somModel.sram_ptr[6][211]=3;
sos_loop[0].somModel.sram_dat[6][212][0]=96'h55b0;
sos_loop[0].somModel.sram_ptr[6][212]=3;
sos_loop[0].somModel.sram_dat[6][213][0]=96'h9ce1;
sos_loop[0].somModel.sram_ptr[6][213]=3;
sos_loop[0].somModel.sram_dat[6][214][0]=96'h981a;
sos_loop[0].somModel.sram_ptr[6][214]=3;
sos_loop[0].somModel.sram_dat[6][215][0]=96'hbc49;
sos_loop[0].somModel.sram_ptr[6][215]=3;
sos_loop[0].somModel.sram_dat[6][216][0]=96'h2f11;
sos_loop[0].somModel.sram_ptr[6][216]=3;
sos_loop[0].somModel.sram_dat[6][217][0]=96'hdfe5;
sos_loop[0].somModel.sram_ptr[6][217]=3;
sos_loop[0].somModel.sram_dat[6][218][0]=96'h261b;
sos_loop[0].somModel.sram_ptr[6][218]=3;
sos_loop[0].somModel.sram_dat[6][219][0]=96'h297f;
sos_loop[0].somModel.sram_ptr[6][219]=3;
sos_loop[0].somModel.sram_dat[6][220][0]=96'h2d7d;
sos_loop[0].somModel.sram_ptr[6][220]=3;
sos_loop[0].somModel.sram_dat[6][221][0]=96'hee8;
sos_loop[0].somModel.sram_ptr[6][221]=3;
sos_loop[0].somModel.sram_dat[6][222][0]=96'h4561;
sos_loop[0].somModel.sram_ptr[6][222]=3;
sos_loop[0].somModel.sram_dat[6][223][0]=96'hc4c2;
sos_loop[0].somModel.sram_ptr[6][223]=3;
sos_loop[0].somModel.sram_dat[6][224][0]=96'ha32d;
sos_loop[0].somModel.sram_ptr[6][224]=3;
sos_loop[0].somModel.sram_dat[6][225][0]=96'hff23;
sos_loop[0].somModel.sram_ptr[6][225]=3;
sos_loop[0].somModel.sram_dat[6][226][0]=96'hd60a;
sos_loop[0].somModel.sram_ptr[6][226]=3;
sos_loop[0].somModel.sram_dat[6][227][0]=96'h7305;
sos_loop[0].somModel.sram_ptr[6][227]=3;
sos_loop[0].somModel.sram_dat[6][228][0]=96'h8bb6;
sos_loop[0].somModel.sram_ptr[6][228]=3;
sos_loop[0].somModel.sram_dat[6][229][0]=96'hac8c;
sos_loop[0].somModel.sram_ptr[6][229]=3;
sos_loop[0].somModel.sram_dat[6][230][0]=96'h8af0;
sos_loop[0].somModel.sram_ptr[6][230]=3;
sos_loop[0].somModel.sram_dat[6][231][0]=96'h7c83;
sos_loop[0].somModel.sram_ptr[6][231]=3;
sos_loop[0].somModel.sram_dat[6][232][0]=96'he1cf;
sos_loop[0].somModel.sram_ptr[6][232]=3;
sos_loop[0].somModel.sram_dat[6][233][0]=96'he86c;
sos_loop[0].somModel.sram_ptr[6][233]=3;
sos_loop[0].somModel.sram_dat[6][234][0]=96'h8c42;
sos_loop[0].somModel.sram_ptr[6][234]=3;
sos_loop[0].somModel.sram_dat[6][235][0]=96'h5f0;
sos_loop[0].somModel.sram_ptr[6][235]=3;
sos_loop[0].somModel.sram_dat[6][236][0]=96'h7074;
sos_loop[0].somModel.sram_ptr[6][236]=3;
sos_loop[0].somModel.sram_dat[6][237][0]=96'h14a6;
sos_loop[0].somModel.sram_ptr[6][237]=3;
sos_loop[0].somModel.sram_dat[6][238][0]=96'h576;
sos_loop[0].somModel.sram_ptr[6][238]=3;
sos_loop[0].somModel.sram_dat[6][239][0]=96'h5b0b;
sos_loop[0].somModel.sram_ptr[6][239]=3;
sos_loop[0].somModel.sram_dat[6][240][0]=96'h4967;
sos_loop[0].somModel.sram_ptr[6][240]=3;
sos_loop[0].somModel.sram_dat[6][241][0]=96'h8e5;
sos_loop[0].somModel.sram_ptr[6][241]=3;
sos_loop[0].somModel.sram_dat[6][242][0]=96'h5734;
sos_loop[0].somModel.sram_ptr[6][242]=3;
sos_loop[0].somModel.sram_dat[6][243][0]=96'h77b3;
sos_loop[0].somModel.sram_ptr[6][243]=3;
sos_loop[0].somModel.sram_dat[6][244][0]=96'hde81;
sos_loop[0].somModel.sram_ptr[6][244]=3;
sos_loop[0].somModel.sram_dat[6][245][0]=96'h9d79;
sos_loop[0].somModel.sram_ptr[6][245]=3;
sos_loop[0].somModel.sram_dat[6][246][0]=96'he3fe;
sos_loop[0].somModel.sram_ptr[6][246]=3;
sos_loop[0].somModel.sram_dat[6][247][0]=96'h4a66;
sos_loop[0].somModel.sram_ptr[6][247]=3;
sos_loop[0].somModel.sram_dat[6][248][0]=96'hcb9e;
sos_loop[0].somModel.sram_ptr[6][248]=3;
sos_loop[0].somModel.sram_dat[6][249][0]=96'hc1e;
sos_loop[0].somModel.sram_ptr[6][249]=3;
sos_loop[0].somModel.sram_dat[6][250][0]=96'hda01;
sos_loop[0].somModel.sram_ptr[6][250]=3;
sos_loop[0].somModel.sram_dat[6][251][0]=96'hfc70;
sos_loop[0].somModel.sram_ptr[6][251]=3;
sos_loop[0].somModel.sram_dat[6][252][0]=96'h35e4;
sos_loop[0].somModel.sram_ptr[6][252]=3;
sos_loop[0].somModel.sram_dat[6][253][0]=96'h1924;
sos_loop[0].somModel.sram_ptr[6][253]=3;
sos_loop[0].somModel.sram_dat[6][254][0]=96'hcb60;
sos_loop[0].somModel.sram_ptr[6][254]=3;
sos_loop[0].somModel.sram_dat[6][255][0]=96'hcb3;
sos_loop[0].somModel.sram_ptr[6][255]=3;
sos_loop[0].somModel.sram_dat[6][256][0]=96'h7107;
sos_loop[0].somModel.sram_ptr[6][256]=3;
sos_loop[0].somModel.sram_dat[6][257][0]=96'hef06;
sos_loop[0].somModel.sram_ptr[6][257]=3;
sos_loop[0].somModel.sram_dat[6][258][0]=96'hb915;
sos_loop[0].somModel.sram_ptr[6][258]=3;
sos_loop[0].somModel.sram_dat[6][259][0]=96'h569e;
sos_loop[0].somModel.sram_ptr[6][259]=3;
sos_loop[0].somModel.sram_dat[6][260][0]=96'ha5c6;
sos_loop[0].somModel.sram_ptr[6][260]=3;
sos_loop[0].somModel.sram_dat[6][261][0]=96'h561;
sos_loop[0].somModel.sram_ptr[6][261]=3;
sos_loop[0].somModel.sram_dat[6][262][0]=96'h543c;
sos_loop[0].somModel.sram_ptr[6][262]=3;
sos_loop[0].somModel.sram_dat[6][263][0]=96'hf887;
sos_loop[0].somModel.sram_ptr[6][263]=3;
sos_loop[0].somModel.sram_dat[6][264][0]=96'h2449;
sos_loop[0].somModel.sram_ptr[6][264]=3;
sos_loop[0].somModel.sram_dat[6][265][0]=96'haa1;
sos_loop[0].somModel.sram_ptr[6][265]=3;
sos_loop[0].somModel.sram_dat[6][266][0]=96'h20fc;
sos_loop[0].somModel.sram_ptr[6][266]=3;
sos_loop[0].somModel.sram_dat[6][267][0]=96'h19c6;
sos_loop[0].somModel.sram_ptr[6][267]=3;
sos_loop[0].somModel.sram_dat[6][268][0]=96'h8d68;
sos_loop[0].somModel.sram_ptr[6][268]=3;
sos_loop[0].somModel.sram_dat[6][269][0]=96'h1fe5;
sos_loop[0].somModel.sram_ptr[6][269]=3;
sos_loop[0].somModel.sram_dat[6][270][0]=96'h8425;
sos_loop[0].somModel.sram_ptr[6][270]=3;
sos_loop[0].somModel.sram_dat[6][271][0]=96'hce2c;
sos_loop[0].somModel.sram_ptr[6][271]=3;
sos_loop[0].somModel.sram_dat[6][272][0]=96'h9e07;
sos_loop[0].somModel.sram_ptr[6][272]=3;
sos_loop[0].somModel.sram_dat[6][273][0]=96'hc360;
sos_loop[0].somModel.sram_ptr[6][273]=3;
sos_loop[0].somModel.sram_dat[6][274][0]=96'h55a6;
sos_loop[0].somModel.sram_ptr[6][274]=3;
sos_loop[0].somModel.sram_dat[6][275][0]=96'hd3ce;
sos_loop[0].somModel.sram_ptr[6][275]=3;
sos_loop[0].somModel.sram_dat[6][276][0]=96'h49ea;
sos_loop[0].somModel.sram_ptr[6][276]=3;
sos_loop[0].somModel.sram_dat[6][277][0]=96'he2e3;
sos_loop[0].somModel.sram_ptr[6][277]=3;
sos_loop[0].somModel.sram_dat[6][278][0]=96'h2b4e;
sos_loop[0].somModel.sram_ptr[6][278]=3;
sos_loop[0].somModel.sram_dat[6][279][0]=96'h8ad9;
sos_loop[0].somModel.sram_ptr[6][279]=3;
sos_loop[0].somModel.sram_dat[6][280][0]=96'h105a;
sos_loop[0].somModel.sram_ptr[6][280]=3;
sos_loop[0].somModel.sram_dat[6][281][0]=96'h279;
sos_loop[0].somModel.sram_ptr[6][281]=3;
sos_loop[0].somModel.sram_dat[6][282][0]=96'h933b;
sos_loop[0].somModel.sram_ptr[6][282]=3;
sos_loop[0].somModel.sram_dat[6][283][0]=96'ha7d8;
sos_loop[0].somModel.sram_ptr[6][283]=3;
sos_loop[0].somModel.sram_dat[6][284][0]=96'h1660;
sos_loop[0].somModel.sram_ptr[6][284]=3;
sos_loop[0].somModel.sram_dat[6][285][0]=96'h2599;
sos_loop[0].somModel.sram_ptr[6][285]=3;
sos_loop[0].somModel.sram_dat[6][286][0]=96'h8360;
sos_loop[0].somModel.sram_ptr[6][286]=3;
sos_loop[0].somModel.sram_dat[6][287][0]=96'h4e54;
sos_loop[0].somModel.sram_ptr[6][287]=3;
sos_loop[0].somModel.sram_dat[6][288][0]=96'h8196;
sos_loop[0].somModel.sram_ptr[6][288]=3;
sos_loop[0].somModel.sram_dat[6][289][0]=96'hc74f;
sos_loop[0].somModel.sram_ptr[6][289]=3;
sos_loop[0].somModel.sram_dat[6][290][0]=96'hdbe6;
sos_loop[0].somModel.sram_ptr[6][290]=3;
sos_loop[0].somModel.sram_dat[6][291][0]=96'hbe67;
sos_loop[0].somModel.sram_ptr[6][291]=3;
sos_loop[0].somModel.sram_dat[6][292][0]=96'h3b66;
sos_loop[0].somModel.sram_ptr[6][292]=3;
sos_loop[0].somModel.sram_dat[6][293][0]=96'hf5d;
sos_loop[0].somModel.sram_ptr[6][293]=3;
sos_loop[0].somModel.sram_dat[6][294][0]=96'h3e97;
sos_loop[0].somModel.sram_ptr[6][294]=3;
sos_loop[0].somModel.sram_dat[6][295][0]=96'h77cb;
sos_loop[0].somModel.sram_ptr[6][295]=3;
sos_loop[0].somModel.sram_dat[6][296][0]=96'h4ffa;
sos_loop[0].somModel.sram_ptr[6][296]=3;
sos_loop[0].somModel.sram_dat[6][297][0]=96'h5a27;
sos_loop[0].somModel.sram_ptr[6][297]=3;
sos_loop[0].somModel.sram_dat[6][298][0]=96'h4f4a;
sos_loop[0].somModel.sram_ptr[6][298]=3;
sos_loop[0].somModel.sram_dat[6][299][0]=96'h89b;
sos_loop[0].somModel.sram_ptr[6][299]=3;
sos_loop[0].somModel.sram_dat[6][300][0]=96'h431f;
sos_loop[0].somModel.sram_ptr[6][300]=3;
sos_loop[0].somModel.sram_dat[6][301][0]=96'hf164;
sos_loop[0].somModel.sram_ptr[6][301]=3;
sos_loop[0].somModel.sram_dat[6][302][0]=96'hae3b;
sos_loop[0].somModel.sram_ptr[6][302]=3;
sos_loop[0].somModel.sram_dat[6][303][0]=96'h4616;
sos_loop[0].somModel.sram_ptr[6][303]=3;
sos_loop[0].somModel.sram_dat[6][304][0]=96'he0cf;
sos_loop[0].somModel.sram_ptr[6][304]=3;
sos_loop[0].somModel.sram_dat[6][305][0]=96'h6917;
sos_loop[0].somModel.sram_ptr[6][305]=3;
sos_loop[0].somModel.sram_dat[6][306][0]=96'h2d00;
sos_loop[0].somModel.sram_ptr[6][306]=3;
sos_loop[0].somModel.sram_dat[6][307][0]=96'h75f9;
sos_loop[0].somModel.sram_ptr[6][307]=3;
sos_loop[0].somModel.sram_dat[6][308][0]=96'h7b29;
sos_loop[0].somModel.sram_ptr[6][308]=3;
sos_loop[0].somModel.sram_dat[6][309][0]=96'h18be;
sos_loop[0].somModel.sram_ptr[6][309]=3;
sos_loop[0].somModel.sram_dat[6][310][0]=96'h87d2;
sos_loop[0].somModel.sram_ptr[6][310]=3;
sos_loop[0].somModel.sram_dat[6][311][0]=96'h3974;
sos_loop[0].somModel.sram_ptr[6][311]=3;
sos_loop[0].somModel.sram_dat[6][312][0]=96'h5c4;
sos_loop[0].somModel.sram_ptr[6][312]=3;
sos_loop[0].somModel.sram_dat[6][313][0]=96'h18b0;
sos_loop[0].somModel.sram_ptr[6][313]=3;
sos_loop[0].somModel.sram_dat[6][314][0]=96'h89fd;
sos_loop[0].somModel.sram_ptr[6][314]=3;
sos_loop[0].somModel.sram_dat[6][315][0]=96'h2c4e;
sos_loop[0].somModel.sram_ptr[6][315]=3;
sos_loop[0].somModel.sram_dat[6][316][0]=96'h417a;
sos_loop[0].somModel.sram_ptr[6][316]=3;
sos_loop[0].somModel.sram_dat[6][317][0]=96'h4888;
sos_loop[0].somModel.sram_ptr[6][317]=3;
sos_loop[0].somModel.sram_dat[6][318][0]=96'h7064;
sos_loop[0].somModel.sram_ptr[6][318]=3;
sos_loop[0].somModel.sram_dat[6][319][0]=96'hb2bf;
sos_loop[0].somModel.sram_ptr[6][319]=3;
sos_loop[0].somModel.sram_dat[6][320][0]=96'h9d55;
sos_loop[0].somModel.sram_ptr[6][320]=3;
sos_loop[0].somModel.sram_dat[6][321][0]=96'hff62;
sos_loop[0].somModel.sram_ptr[6][321]=3;
sos_loop[0].somModel.sram_dat[6][322][0]=96'hb397;
sos_loop[0].somModel.sram_ptr[6][322]=3;
sos_loop[0].somModel.sram_dat[6][323][0]=96'hbbdd;
sos_loop[0].somModel.sram_ptr[6][323]=3;
sos_loop[0].somModel.sram_dat[6][324][0]=96'h871d;
sos_loop[0].somModel.sram_ptr[6][324]=3;
sos_loop[0].somModel.sram_dat[6][325][0]=96'h6fe6;
sos_loop[0].somModel.sram_ptr[6][325]=3;
sos_loop[0].somModel.sram_dat[6][326][0]=96'hb4f0;
sos_loop[0].somModel.sram_ptr[6][326]=3;
sos_loop[0].somModel.sram_dat[6][327][0]=96'h343b;
sos_loop[0].somModel.sram_ptr[6][327]=3;
sos_loop[0].somModel.sram_dat[6][328][0]=96'h7848;
sos_loop[0].somModel.sram_ptr[6][328]=3;
sos_loop[0].somModel.sram_dat[6][329][0]=96'h826c;
sos_loop[0].somModel.sram_ptr[6][329]=3;
sos_loop[0].somModel.sram_dat[6][330][0]=96'h466e;
sos_loop[0].somModel.sram_ptr[6][330]=3;
sos_loop[0].somModel.sram_dat[6][331][0]=96'h6d50;
sos_loop[0].somModel.sram_ptr[6][331]=3;
sos_loop[0].somModel.sram_dat[6][332][0]=96'h892d;
sos_loop[0].somModel.sram_ptr[6][332]=3;
sos_loop[0].somModel.sram_dat[6][333][0]=96'h8567;
sos_loop[0].somModel.sram_ptr[6][333]=3;
sos_loop[0].somModel.sram_dat[6][334][0]=96'hb0d3;
sos_loop[0].somModel.sram_ptr[6][334]=3;
sos_loop[0].somModel.sram_dat[6][335][0]=96'hc89f;
sos_loop[0].somModel.sram_ptr[6][335]=3;
sos_loop[0].somModel.sram_dat[6][336][0]=96'h2ac3;
sos_loop[0].somModel.sram_ptr[6][336]=3;
sos_loop[0].somModel.sram_dat[6][337][0]=96'h7e5e;
sos_loop[0].somModel.sram_ptr[6][337]=3;
sos_loop[0].somModel.sram_dat[6][338][0]=96'hd4e5;
sos_loop[0].somModel.sram_ptr[6][338]=3;
sos_loop[0].somModel.sram_dat[6][339][0]=96'hd1f0;
sos_loop[0].somModel.sram_ptr[6][339]=3;
sos_loop[0].somModel.sram_dat[6][340][0]=96'h81b0;
sos_loop[0].somModel.sram_ptr[6][340]=3;
sos_loop[0].somModel.sram_dat[6][341][0]=96'hfcdf;
sos_loop[0].somModel.sram_ptr[6][341]=3;
sos_loop[0].somModel.sram_dat[6][342][0]=96'h56e8;
sos_loop[0].somModel.sram_ptr[6][342]=3;
sos_loop[0].somModel.sram_dat[6][343][0]=96'h9ba4;
sos_loop[0].somModel.sram_ptr[6][343]=3;
sos_loop[0].somModel.sram_dat[6][344][0]=96'h9667;
sos_loop[0].somModel.sram_ptr[6][344]=3;
sos_loop[0].somModel.sram_dat[6][345][0]=96'h3024;
sos_loop[0].somModel.sram_ptr[6][345]=3;
sos_loop[0].somModel.sram_dat[6][346][0]=96'he58;
sos_loop[0].somModel.sram_ptr[6][346]=3;
sos_loop[0].somModel.sram_dat[6][347][0]=96'hd571;
sos_loop[0].somModel.sram_ptr[6][347]=3;
sos_loop[0].somModel.sram_dat[6][348][0]=96'h7454;
sos_loop[0].somModel.sram_ptr[6][348]=3;
sos_loop[0].somModel.sram_dat[6][349][0]=96'h11fb;
sos_loop[0].somModel.sram_ptr[6][349]=3;
sos_loop[0].somModel.sram_dat[6][350][0]=96'h6209;
sos_loop[0].somModel.sram_ptr[6][350]=3;
sos_loop[0].somModel.sram_dat[6][351][0]=96'he475;
sos_loop[0].somModel.sram_ptr[6][351]=3;
sos_loop[0].somModel.sram_dat[6][352][0]=96'hc860;
sos_loop[0].somModel.sram_ptr[6][352]=3;
sos_loop[0].somModel.sram_dat[6][353][0]=96'h781;
sos_loop[0].somModel.sram_ptr[6][353]=3;
sos_loop[0].somModel.sram_dat[6][354][0]=96'h2590;
sos_loop[0].somModel.sram_ptr[6][354]=3;
sos_loop[0].somModel.sram_dat[6][355][0]=96'hfa8e;
sos_loop[0].somModel.sram_ptr[6][355]=3;
sos_loop[0].somModel.sram_dat[6][356][0]=96'h3f7d;
sos_loop[0].somModel.sram_ptr[6][356]=3;
sos_loop[0].somModel.sram_dat[6][357][0]=96'h515;
sos_loop[0].somModel.sram_ptr[6][357]=3;
sos_loop[0].somModel.sram_dat[6][358][0]=96'hb9b3;
sos_loop[0].somModel.sram_ptr[6][358]=3;
sos_loop[0].somModel.sram_dat[6][359][0]=96'h6db1;
sos_loop[0].somModel.sram_ptr[6][359]=3;
sos_loop[0].somModel.sram_dat[6][360][0]=96'hcde4;
sos_loop[0].somModel.sram_ptr[6][360]=3;
sos_loop[0].somModel.sram_dat[6][361][0]=96'hce02;
sos_loop[0].somModel.sram_ptr[6][361]=3;
sos_loop[0].somModel.sram_dat[6][362][0]=96'h4a3c;
sos_loop[0].somModel.sram_ptr[6][362]=3;
sos_loop[0].somModel.sram_dat[6][363][0]=96'h8440;
sos_loop[0].somModel.sram_ptr[6][363]=3;
sos_loop[0].somModel.sram_dat[6][364][0]=96'h82a7;
sos_loop[0].somModel.sram_ptr[6][364]=3;
sos_loop[0].somModel.sram_dat[6][365][0]=96'he481;
sos_loop[0].somModel.sram_ptr[6][365]=3;
sos_loop[0].somModel.sram_dat[6][366][0]=96'h1c1b;
sos_loop[0].somModel.sram_ptr[6][366]=3;
sos_loop[0].somModel.sram_dat[6][367][0]=96'h819b;
sos_loop[0].somModel.sram_ptr[6][367]=3;
sos_loop[0].somModel.sram_dat[6][368][0]=96'he56e;
sos_loop[0].somModel.sram_ptr[6][368]=3;
sos_loop[0].somModel.sram_dat[6][369][0]=96'h84c7;
sos_loop[0].somModel.sram_ptr[6][369]=3;
sos_loop[0].somModel.sram_dat[6][370][0]=96'h2c16;
sos_loop[0].somModel.sram_ptr[6][370]=3;
sos_loop[0].somModel.sram_dat[6][371][0]=96'h4fb9;
sos_loop[0].somModel.sram_ptr[6][371]=3;
sos_loop[0].somModel.sram_dat[6][372][0]=96'h5dad;
sos_loop[0].somModel.sram_ptr[6][372]=3;
sos_loop[0].somModel.sram_dat[6][373][0]=96'h4e74;
sos_loop[0].somModel.sram_ptr[6][373]=3;
sos_loop[0].somModel.sram_dat[6][374][0]=96'h30d5;
sos_loop[0].somModel.sram_ptr[6][374]=3;
sos_loop[0].somModel.sram_dat[6][375][0]=96'h41fa;
sos_loop[0].somModel.sram_ptr[6][375]=3;
sos_loop[0].somModel.sram_dat[6][376][0]=96'hbf53;
sos_loop[0].somModel.sram_ptr[6][376]=3;
sos_loop[0].somModel.sram_dat[6][377][0]=96'h901d;
sos_loop[0].somModel.sram_ptr[6][377]=3;
sos_loop[0].somModel.sram_dat[6][378][0]=96'hf3ee;
sos_loop[0].somModel.sram_ptr[6][378]=3;
sos_loop[0].somModel.sram_dat[6][379][0]=96'h9197;
sos_loop[0].somModel.sram_ptr[6][379]=3;
sos_loop[0].somModel.sram_dat[6][380][0]=96'h1aac;
sos_loop[0].somModel.sram_ptr[6][380]=3;
sos_loop[0].somModel.sram_dat[6][381][0]=96'hcc69;
sos_loop[0].somModel.sram_ptr[6][381]=3;
sos_loop[0].somModel.sram_dat[6][382][0]=96'h3722;
sos_loop[0].somModel.sram_ptr[6][382]=3;
sos_loop[0].somModel.sram_dat[6][383][0]=96'hda62;
sos_loop[0].somModel.sram_ptr[6][383]=3;
sos_loop[0].somModel.sram_dat[6][384][0]=96'hc7f6;
sos_loop[0].somModel.sram_ptr[6][384]=3;
sos_loop[0].somModel.sram_dat[6][385][0]=96'he590;
sos_loop[0].somModel.sram_ptr[6][385]=3;
sos_loop[0].somModel.sram_dat[6][386][0]=96'h8354;
sos_loop[0].somModel.sram_ptr[6][386]=3;
sos_loop[0].somModel.sram_dat[6][387][0]=96'hdee4;
sos_loop[0].somModel.sram_ptr[6][387]=3;
sos_loop[0].somModel.sram_dat[6][388][0]=96'h8a42;
sos_loop[0].somModel.sram_ptr[6][388]=3;
sos_loop[0].somModel.sram_dat[6][389][0]=96'h8249;
sos_loop[0].somModel.sram_ptr[6][389]=3;
sos_loop[0].somModel.sram_dat[6][390][0]=96'hd7b2;
sos_loop[0].somModel.sram_ptr[6][390]=3;
sos_loop[0].somModel.sram_dat[6][391][0]=96'hdb8d;
sos_loop[0].somModel.sram_ptr[6][391]=3;
sos_loop[0].somModel.sram_dat[6][392][0]=96'h7dca;
sos_loop[0].somModel.sram_ptr[6][392]=3;
sos_loop[0].somModel.sram_dat[6][393][0]=96'h4cb3;
sos_loop[0].somModel.sram_ptr[6][393]=3;
sos_loop[0].somModel.sram_dat[6][394][0]=96'h7648;
sos_loop[0].somModel.sram_ptr[6][394]=3;
sos_loop[0].somModel.sram_dat[6][395][0]=96'h51a0;
sos_loop[0].somModel.sram_ptr[6][395]=3;
sos_loop[0].somModel.sram_dat[6][396][0]=96'hfce6;
sos_loop[0].somModel.sram_ptr[6][396]=3;
sos_loop[0].somModel.sram_dat[6][397][0]=96'h1a6e;
sos_loop[0].somModel.sram_ptr[6][397]=3;
sos_loop[0].somModel.sram_dat[6][398][0]=96'h4fab;
sos_loop[0].somModel.sram_ptr[6][398]=3;
sos_loop[0].somModel.sram_dat[6][399][0]=96'hb664;
sos_loop[0].somModel.sram_ptr[6][399]=3;
sos_loop[0].somModel.sram_dat[6][400][0]=96'h7466;
sos_loop[0].somModel.sram_ptr[6][400]=3;
sos_loop[0].somModel.sram_dat[6][401][0]=96'h5d91;
sos_loop[0].somModel.sram_ptr[6][401]=3;
sos_loop[0].somModel.sram_dat[6][402][0]=96'ha6d9;
sos_loop[0].somModel.sram_ptr[6][402]=3;
sos_loop[0].somModel.sram_dat[6][403][0]=96'h66a;
sos_loop[0].somModel.sram_ptr[6][403]=3;
sos_loop[0].somModel.sram_dat[6][404][0]=96'h6c8b;
sos_loop[0].somModel.sram_ptr[6][404]=3;
sos_loop[0].somModel.sram_dat[6][405][0]=96'h7561;
sos_loop[0].somModel.sram_ptr[6][405]=3;
sos_loop[0].somModel.sram_dat[6][406][0]=96'h2b5e;
sos_loop[0].somModel.sram_ptr[6][406]=3;
sos_loop[0].somModel.sram_dat[6][407][0]=96'h5f68;
sos_loop[0].somModel.sram_ptr[6][407]=3;
sos_loop[0].somModel.sram_dat[6][408][0]=96'h8d5a;
sos_loop[0].somModel.sram_ptr[6][408]=3;
sos_loop[0].somModel.sram_dat[6][409][0]=96'h5ff9;
sos_loop[0].somModel.sram_ptr[6][409]=3;
sos_loop[0].somModel.sram_dat[6][410][0]=96'haa4a;
sos_loop[0].somModel.sram_ptr[6][410]=3;
sos_loop[0].somModel.sram_dat[6][411][0]=96'h9b48;
sos_loop[0].somModel.sram_ptr[6][411]=3;
sos_loop[0].somModel.sram_dat[6][412][0]=96'hbab5;
sos_loop[0].somModel.sram_ptr[6][412]=3;
sos_loop[0].somModel.sram_dat[6][413][0]=96'he87e;
sos_loop[0].somModel.sram_ptr[6][413]=3;
sos_loop[0].somModel.sram_dat[6][414][0]=96'h27ff;
sos_loop[0].somModel.sram_ptr[6][414]=3;
sos_loop[0].somModel.sram_dat[6][415][0]=96'hdb49;
sos_loop[0].somModel.sram_ptr[6][415]=3;
sos_loop[0].somModel.sram_dat[6][416][0]=96'ha716;
sos_loop[0].somModel.sram_ptr[6][416]=3;
sos_loop[0].somModel.sram_dat[6][417][0]=96'hea5e;
sos_loop[0].somModel.sram_ptr[6][417]=3;
sos_loop[0].somModel.sram_dat[6][418][0]=96'h9813;
sos_loop[0].somModel.sram_ptr[6][418]=3;
sos_loop[0].somModel.sram_dat[6][419][0]=96'h1c2b;
sos_loop[0].somModel.sram_ptr[6][419]=3;
sos_loop[0].somModel.sram_dat[6][420][0]=96'h5490;
sos_loop[0].somModel.sram_ptr[6][420]=3;
sos_loop[0].somModel.sram_dat[6][421][0]=96'hdbbc;
sos_loop[0].somModel.sram_ptr[6][421]=3;
sos_loop[0].somModel.sram_dat[6][422][0]=96'hba73;
sos_loop[0].somModel.sram_ptr[6][422]=3;
sos_loop[0].somModel.sram_dat[6][423][0]=96'h22b8;
sos_loop[0].somModel.sram_ptr[6][423]=3;
sos_loop[0].somModel.sram_dat[6][424][0]=96'h4004;
sos_loop[0].somModel.sram_ptr[6][424]=3;
sos_loop[0].somModel.sram_dat[6][425][0]=96'h1d02;
sos_loop[0].somModel.sram_ptr[6][425]=3;
sos_loop[0].somModel.sram_dat[6][426][0]=96'h32bd;
sos_loop[0].somModel.sram_ptr[6][426]=3;
sos_loop[0].somModel.sram_dat[6][427][0]=96'h5a87;
sos_loop[0].somModel.sram_ptr[6][427]=3;
sos_loop[0].somModel.sram_dat[6][428][0]=96'h1835;
sos_loop[0].somModel.sram_ptr[6][428]=3;
sos_loop[0].somModel.sram_dat[6][429][0]=96'h348;
sos_loop[0].somModel.sram_ptr[6][429]=3;
sos_loop[0].somModel.sram_dat[6][430][0]=96'h7db8;
sos_loop[0].somModel.sram_ptr[6][430]=3;
sos_loop[0].somModel.sram_dat[6][431][0]=96'h53a0;
sos_loop[0].somModel.sram_ptr[6][431]=3;
sos_loop[0].somModel.sram_dat[6][432][0]=96'h94a;
sos_loop[0].somModel.sram_ptr[6][432]=3;
sos_loop[0].somModel.sram_dat[6][433][0]=96'h68a9;
sos_loop[0].somModel.sram_ptr[6][433]=3;
sos_loop[0].somModel.sram_dat[6][434][0]=96'h6588;
sos_loop[0].somModel.sram_ptr[6][434]=3;
sos_loop[0].somModel.sram_dat[6][435][0]=96'h54d3;
sos_loop[0].somModel.sram_ptr[6][435]=3;
sos_loop[0].somModel.sram_dat[6][436][0]=96'h7b1e;
sos_loop[0].somModel.sram_ptr[6][436]=3;
sos_loop[0].somModel.sram_dat[6][437][0]=96'h6a07;
sos_loop[0].somModel.sram_ptr[6][437]=3;
sos_loop[0].somModel.sram_dat[6][438][0]=96'hecf4;
sos_loop[0].somModel.sram_ptr[6][438]=3;
sos_loop[0].somModel.sram_dat[6][439][0]=96'h75f1;
sos_loop[0].somModel.sram_ptr[6][439]=3;
sos_loop[0].somModel.sram_dat[6][440][0]=96'h17b4;
sos_loop[0].somModel.sram_ptr[6][440]=3;
sos_loop[0].somModel.sram_dat[6][441][0]=96'h8fcf;
sos_loop[0].somModel.sram_ptr[6][441]=3;
sos_loop[0].somModel.sram_dat[6][442][0]=96'hfd38;
sos_loop[0].somModel.sram_ptr[6][442]=3;
sos_loop[0].somModel.sram_dat[6][443][0]=96'h2d2;
sos_loop[0].somModel.sram_ptr[6][443]=3;
sos_loop[0].somModel.sram_dat[6][444][0]=96'hc881;
sos_loop[0].somModel.sram_ptr[6][444]=3;
sos_loop[0].somModel.sram_dat[6][445][0]=96'hbb36;
sos_loop[0].somModel.sram_ptr[6][445]=3;
sos_loop[0].somModel.sram_dat[6][446][0]=96'h86ff;
sos_loop[0].somModel.sram_ptr[6][446]=3;
sos_loop[0].somModel.sram_dat[6][447][0]=96'ha23f;
sos_loop[0].somModel.sram_ptr[6][447]=3;
sos_loop[0].somModel.sram_dat[6][448][0]=96'hd8ec;
sos_loop[0].somModel.sram_ptr[6][448]=3;
sos_loop[0].somModel.sram_dat[6][449][0]=96'h5f93;
sos_loop[0].somModel.sram_ptr[6][449]=3;
sos_loop[0].somModel.sram_dat[6][450][0]=96'hbc1;
sos_loop[0].somModel.sram_ptr[6][450]=3;
sos_loop[0].somModel.sram_dat[6][451][0]=96'h144;
sos_loop[0].somModel.sram_ptr[6][451]=3;
sos_loop[0].somModel.sram_dat[6][452][0]=96'hfdbe;
sos_loop[0].somModel.sram_ptr[6][452]=3;
sos_loop[0].somModel.sram_dat[6][453][0]=96'h70f4;
sos_loop[0].somModel.sram_ptr[6][453]=3;
sos_loop[0].somModel.sram_dat[6][454][0]=96'h5006;
sos_loop[0].somModel.sram_ptr[6][454]=3;
sos_loop[0].somModel.sram_dat[6][455][0]=96'h4772;
sos_loop[0].somModel.sram_ptr[6][455]=3;
sos_loop[0].somModel.sram_dat[6][456][0]=96'h1aa8;
sos_loop[0].somModel.sram_ptr[6][456]=3;
sos_loop[0].somModel.sram_dat[6][457][0]=96'hdd72;
sos_loop[0].somModel.sram_ptr[6][457]=3;
sos_loop[0].somModel.sram_dat[6][458][0]=96'h2ec4;
sos_loop[0].somModel.sram_ptr[6][458]=3;
sos_loop[0].somModel.sram_dat[6][459][0]=96'h33f9;
sos_loop[0].somModel.sram_ptr[6][459]=3;
sos_loop[0].somModel.sram_dat[6][460][0]=96'ha3f3;
sos_loop[0].somModel.sram_ptr[6][460]=3;
sos_loop[0].somModel.sram_dat[6][461][0]=96'h8144;
sos_loop[0].somModel.sram_ptr[6][461]=3;
sos_loop[0].somModel.sram_dat[6][462][0]=96'h6971;
sos_loop[0].somModel.sram_ptr[6][462]=3;
sos_loop[0].somModel.sram_dat[6][463][0]=96'h3a0f;
sos_loop[0].somModel.sram_ptr[6][463]=3;
sos_loop[0].somModel.sram_dat[6][464][0]=96'hf3b3;
sos_loop[0].somModel.sram_ptr[6][464]=3;
sos_loop[0].somModel.sram_dat[6][465][0]=96'h4c3;
sos_loop[0].somModel.sram_ptr[6][465]=3;
sos_loop[0].somModel.sram_dat[6][466][0]=96'h97a2;
sos_loop[0].somModel.sram_ptr[6][466]=3;
sos_loop[0].somModel.sram_dat[6][467][0]=96'h191e;
sos_loop[0].somModel.sram_ptr[6][467]=3;
sos_loop[0].somModel.sram_dat[6][468][0]=96'h4c9d;
sos_loop[0].somModel.sram_ptr[6][468]=3;
sos_loop[0].somModel.sram_dat[6][469][0]=96'h1c56;
sos_loop[0].somModel.sram_ptr[6][469]=3;
sos_loop[0].somModel.sram_dat[6][470][0]=96'h4f2e;
sos_loop[0].somModel.sram_ptr[6][470]=3;
sos_loop[0].somModel.sram_dat[6][471][0]=96'h7a32;
sos_loop[0].somModel.sram_ptr[6][471]=3;
sos_loop[0].somModel.sram_dat[6][472][0]=96'he58e;
sos_loop[0].somModel.sram_ptr[6][472]=3;
sos_loop[0].somModel.sram_dat[6][473][0]=96'hfc5;
sos_loop[0].somModel.sram_ptr[6][473]=3;
sos_loop[0].somModel.sram_dat[6][474][0]=96'h30ab;
sos_loop[0].somModel.sram_ptr[6][474]=3;
sos_loop[0].somModel.sram_dat[6][475][0]=96'h8377;
sos_loop[0].somModel.sram_ptr[6][475]=3;
sos_loop[0].somModel.sram_dat[6][476][0]=96'hd368;
sos_loop[0].somModel.sram_ptr[6][476]=3;
sos_loop[0].somModel.sram_dat[6][477][0]=96'h6d1d;
sos_loop[0].somModel.sram_ptr[6][477]=3;
sos_loop[0].somModel.sram_dat[6][478][0]=96'h23a3;
sos_loop[0].somModel.sram_ptr[6][478]=3;
sos_loop[0].somModel.sram_dat[6][479][0]=96'h4845;
sos_loop[0].somModel.sram_ptr[6][479]=3;
sos_loop[0].somModel.sram_dat[6][480][0]=96'h992e;
sos_loop[0].somModel.sram_ptr[6][480]=3;
sos_loop[0].somModel.sram_dat[6][481][0]=96'h9aad;
sos_loop[0].somModel.sram_ptr[6][481]=3;
sos_loop[0].somModel.sram_dat[6][482][0]=96'hc17;
sos_loop[0].somModel.sram_ptr[6][482]=3;
sos_loop[0].somModel.sram_dat[6][483][0]=96'hce74;
sos_loop[0].somModel.sram_ptr[6][483]=3;
sos_loop[0].somModel.sram_dat[6][484][0]=96'ha3bc;
sos_loop[0].somModel.sram_ptr[6][484]=3;
sos_loop[0].somModel.sram_dat[6][485][0]=96'haf3e;
sos_loop[0].somModel.sram_ptr[6][485]=3;
sos_loop[0].somModel.sram_dat[6][486][0]=96'hf44a;
sos_loop[0].somModel.sram_ptr[6][486]=3;
sos_loop[0].somModel.sram_dat[6][487][0]=96'habdc;
sos_loop[0].somModel.sram_ptr[6][487]=3;
sos_loop[0].somModel.sram_dat[6][488][0]=96'h1ffa;
sos_loop[0].somModel.sram_ptr[6][488]=3;
sos_loop[0].somModel.sram_dat[6][489][0]=96'hbbe8;
sos_loop[0].somModel.sram_ptr[6][489]=3;
sos_loop[0].somModel.sram_dat[6][490][0]=96'hce02;
sos_loop[0].somModel.sram_ptr[6][490]=3;
sos_loop[0].somModel.sram_dat[6][491][0]=96'hf7a;
sos_loop[0].somModel.sram_ptr[6][491]=3;
sos_loop[0].somModel.sram_dat[6][492][0]=96'hb92;
sos_loop[0].somModel.sram_ptr[6][492]=3;
sos_loop[0].somModel.sram_dat[6][493][0]=96'h371a;
sos_loop[0].somModel.sram_ptr[6][493]=3;
sos_loop[0].somModel.sram_dat[6][494][0]=96'h5154;
sos_loop[0].somModel.sram_ptr[6][494]=3;
sos_loop[0].somModel.sram_dat[6][495][0]=96'h244d;
sos_loop[0].somModel.sram_ptr[6][495]=3;
sos_loop[0].somModel.sram_dat[6][496][0]=96'hd841;
sos_loop[0].somModel.sram_ptr[6][496]=3;
sos_loop[0].somModel.sram_dat[6][497][0]=96'h7799;
sos_loop[0].somModel.sram_ptr[6][497]=3;
sos_loop[0].somModel.sram_dat[6][498][0]=96'h4853;
sos_loop[0].somModel.sram_ptr[6][498]=3;
sos_loop[0].somModel.sram_dat[6][499][0]=96'h9615;
sos_loop[0].somModel.sram_ptr[6][499]=3;
sos_loop[0].somModel.sram_dat[6][500][0]=96'h25af;
sos_loop[0].somModel.sram_ptr[6][500]=3;
sos_loop[0].somModel.sram_dat[6][501][0]=96'h25f9;
sos_loop[0].somModel.sram_ptr[6][501]=3;
sos_loop[0].somModel.sram_dat[6][502][0]=96'h2c36;
sos_loop[0].somModel.sram_ptr[6][502]=3;
sos_loop[0].somModel.sram_dat[6][503][0]=96'h6575;
sos_loop[0].somModel.sram_ptr[6][503]=3;
sos_loop[0].somModel.sram_dat[6][504][0]=96'h3684;
sos_loop[0].somModel.sram_ptr[6][504]=3;
sos_loop[0].somModel.sram_dat[6][505][0]=96'hf639;
sos_loop[0].somModel.sram_ptr[6][505]=3;
sos_loop[0].somModel.sram_dat[6][506][0]=96'h26d1;
sos_loop[0].somModel.sram_ptr[6][506]=3;
sos_loop[0].somModel.sram_dat[6][507][0]=96'h13dd;
sos_loop[0].somModel.sram_ptr[6][507]=3;
sos_loop[0].somModel.sram_dat[6][508][0]=96'h3335;
sos_loop[0].somModel.sram_ptr[6][508]=3;
sos_loop[0].somModel.sram_dat[6][509][0]=96'he6ea;
sos_loop[0].somModel.sram_ptr[6][509]=3;
sos_loop[0].somModel.sram_dat[6][510][0]=96'h1403;
sos_loop[0].somModel.sram_ptr[6][510]=3;
sos_loop[0].somModel.sram_dat[6][511][0]=96'hb48a;
sos_loop[0].somModel.sram_ptr[6][511]=3;
sos_loop[0].somModel.sram_dat[6][512][0]=96'h3a1b;
sos_loop[0].somModel.sram_ptr[6][512]=3;
sos_loop[0].somModel.sram_dat[6][513][0]=96'hc0f4;
sos_loop[0].somModel.sram_ptr[6][513]=3;
sos_loop[0].somModel.sram_dat[6][514][0]=96'hb6f5;
sos_loop[0].somModel.sram_ptr[6][514]=3;
sos_loop[0].somModel.sram_dat[6][515][0]=96'h5c2f;
sos_loop[0].somModel.sram_ptr[6][515]=3;
sos_loop[0].somModel.sram_dat[6][516][0]=96'h62e1;
sos_loop[0].somModel.sram_ptr[6][516]=3;
sos_loop[0].somModel.sram_dat[6][517][0]=96'hc121;
sos_loop[0].somModel.sram_ptr[6][517]=3;
sos_loop[0].somModel.sram_dat[6][518][0]=96'hc629;
sos_loop[0].somModel.sram_ptr[6][518]=3;
sos_loop[0].somModel.sram_dat[6][519][0]=96'h19d2;
sos_loop[0].somModel.sram_ptr[6][519]=3;
sos_loop[0].somModel.sram_dat[6][520][0]=96'h9600;
sos_loop[0].somModel.sram_ptr[6][520]=3;
sos_loop[0].somModel.sram_dat[6][521][0]=96'hb54;
sos_loop[0].somModel.sram_ptr[6][521]=3;
sos_loop[0].somModel.sram_dat[6][522][0]=96'hd9db;
sos_loop[0].somModel.sram_ptr[6][522]=3;
sos_loop[0].somModel.sram_dat[6][523][0]=96'h284a;
sos_loop[0].somModel.sram_ptr[6][523]=3;
sos_loop[0].somModel.sram_dat[6][524][0]=96'h6511;
sos_loop[0].somModel.sram_ptr[6][524]=3;
sos_loop[0].somModel.sram_dat[6][525][0]=96'hb42e;
sos_loop[0].somModel.sram_ptr[6][525]=3;
sos_loop[0].somModel.sram_dat[6][526][0]=96'ha05a;
sos_loop[0].somModel.sram_ptr[6][526]=3;
sos_loop[0].somModel.sram_dat[6][527][0]=96'h4f13;
sos_loop[0].somModel.sram_ptr[6][527]=3;
sos_loop[0].somModel.sram_dat[6][528][0]=96'h5ae;
sos_loop[0].somModel.sram_ptr[6][528]=3;
sos_loop[0].somModel.sram_dat[6][529][0]=96'h2d8c;
sos_loop[0].somModel.sram_ptr[6][529]=3;
sos_loop[0].somModel.sram_dat[6][530][0]=96'h2bff;
sos_loop[0].somModel.sram_ptr[6][530]=3;
sos_loop[0].somModel.sram_dat[6][531][0]=96'h9abe;
sos_loop[0].somModel.sram_ptr[6][531]=3;
sos_loop[0].somModel.sram_dat[6][532][0]=96'hcfd9;
sos_loop[0].somModel.sram_ptr[6][532]=3;
sos_loop[0].somModel.sram_dat[6][533][0]=96'h3957;
sos_loop[0].somModel.sram_ptr[6][533]=3;
sos_loop[0].somModel.sram_dat[6][534][0]=96'h4efb;
sos_loop[0].somModel.sram_ptr[6][534]=3;
sos_loop[0].somModel.sram_dat[6][535][0]=96'hdd5e;
sos_loop[0].somModel.sram_ptr[6][535]=3;
sos_loop[0].somModel.sram_dat[6][536][0]=96'h800e;
sos_loop[0].somModel.sram_ptr[6][536]=3;
sos_loop[0].somModel.sram_dat[6][537][0]=96'h1697;
sos_loop[0].somModel.sram_ptr[6][537]=3;
sos_loop[0].somModel.sram_dat[6][538][0]=96'h42ce;
sos_loop[0].somModel.sram_ptr[6][538]=3;
sos_loop[0].somModel.sram_dat[6][539][0]=96'hbcbf;
sos_loop[0].somModel.sram_ptr[6][539]=3;
sos_loop[0].somModel.sram_dat[6][540][0]=96'h8541;
sos_loop[0].somModel.sram_ptr[6][540]=3;
sos_loop[0].somModel.sram_dat[6][541][0]=96'h85d1;
sos_loop[0].somModel.sram_ptr[6][541]=3;
sos_loop[0].somModel.sram_dat[6][542][0]=96'h3385;
sos_loop[0].somModel.sram_ptr[6][542]=3;
sos_loop[0].somModel.sram_dat[6][543][0]=96'h708c;
sos_loop[0].somModel.sram_ptr[6][543]=3;
sos_loop[0].somModel.sram_dat[6][544][0]=96'h2082;
sos_loop[0].somModel.sram_ptr[6][544]=3;
sos_loop[0].somModel.sram_dat[6][545][0]=96'h55b;
sos_loop[0].somModel.sram_ptr[6][545]=3;
sos_loop[0].somModel.sram_dat[6][546][0]=96'h15db;
sos_loop[0].somModel.sram_ptr[6][546]=3;
sos_loop[0].somModel.sram_dat[6][547][0]=96'h614f;
sos_loop[0].somModel.sram_ptr[6][547]=3;
sos_loop[0].somModel.sram_dat[6][548][0]=96'h13b4;
sos_loop[0].somModel.sram_ptr[6][548]=3;
sos_loop[0].somModel.sram_dat[6][549][0]=96'h4a8b;
sos_loop[0].somModel.sram_ptr[6][549]=3;
sos_loop[0].somModel.sram_dat[6][550][0]=96'hd328;
sos_loop[0].somModel.sram_ptr[6][550]=3;
sos_loop[0].somModel.sram_dat[6][551][0]=96'h2219;
sos_loop[0].somModel.sram_ptr[6][551]=3;
sos_loop[0].somModel.sram_dat[6][552][0]=96'hfdef;
sos_loop[0].somModel.sram_ptr[6][552]=3;
sos_loop[0].somModel.sram_dat[6][553][0]=96'hcab1;
sos_loop[0].somModel.sram_ptr[6][553]=3;
sos_loop[0].somModel.sram_dat[6][554][0]=96'h8dc9;
sos_loop[0].somModel.sram_ptr[6][554]=3;
sos_loop[0].somModel.sram_dat[6][555][0]=96'h8a3e;
sos_loop[0].somModel.sram_ptr[6][555]=3;
sos_loop[0].somModel.sram_dat[6][556][0]=96'h2949;
sos_loop[0].somModel.sram_ptr[6][556]=3;
sos_loop[0].somModel.sram_dat[6][557][0]=96'hd515;
sos_loop[0].somModel.sram_ptr[6][557]=3;
sos_loop[0].somModel.sram_dat[6][558][0]=96'ha7ab;
sos_loop[0].somModel.sram_ptr[6][558]=3;
sos_loop[0].somModel.sram_dat[6][559][0]=96'h8155;
sos_loop[0].somModel.sram_ptr[6][559]=3;
sos_loop[0].somModel.sram_dat[6][560][0]=96'hbbc5;
sos_loop[0].somModel.sram_ptr[6][560]=3;
sos_loop[0].somModel.sram_dat[6][561][0]=96'h5035;
sos_loop[0].somModel.sram_ptr[6][561]=3;
sos_loop[0].somModel.sram_dat[6][562][0]=96'hb93f;
sos_loop[0].somModel.sram_ptr[6][562]=3;
sos_loop[0].somModel.sram_dat[6][563][0]=96'h37bb;
sos_loop[0].somModel.sram_ptr[6][563]=3;
sos_loop[0].somModel.sram_dat[6][564][0]=96'h6387;
sos_loop[0].somModel.sram_ptr[6][564]=3;
sos_loop[0].somModel.sram_dat[6][565][0]=96'h338f;
sos_loop[0].somModel.sram_ptr[6][565]=3;
sos_loop[0].somModel.sram_dat[6][566][0]=96'h26a6;
sos_loop[0].somModel.sram_ptr[6][566]=3;
sos_loop[0].somModel.sram_dat[6][567][0]=96'h206d;
sos_loop[0].somModel.sram_ptr[6][567]=3;
sos_loop[0].somModel.sram_dat[6][568][0]=96'h8535;
sos_loop[0].somModel.sram_ptr[6][568]=3;
sos_loop[0].somModel.sram_dat[6][569][0]=96'h1b88;
sos_loop[0].somModel.sram_ptr[6][569]=3;
sos_loop[0].somModel.sram_dat[6][570][0]=96'hfbe6;
sos_loop[0].somModel.sram_ptr[6][570]=3;
sos_loop[0].somModel.sram_dat[6][571][0]=96'he4bf;
sos_loop[0].somModel.sram_ptr[6][571]=3;
sos_loop[0].somModel.sram_dat[6][572][0]=96'ha5a6;
sos_loop[0].somModel.sram_ptr[6][572]=3;
sos_loop[0].somModel.sram_dat[6][573][0]=96'h9f00;
sos_loop[0].somModel.sram_ptr[6][573]=3;
sos_loop[0].somModel.sram_dat[6][574][0]=96'h6530;
sos_loop[0].somModel.sram_ptr[6][574]=3;
sos_loop[0].somModel.sram_dat[6][575][0]=96'h37d5;
sos_loop[0].somModel.sram_ptr[6][575]=3;
sos_loop[0].somModel.sram_dat[6][576][0]=96'h9b09;
sos_loop[0].somModel.sram_ptr[6][576]=3;
sos_loop[0].somModel.sram_dat[6][577][0]=96'ha8bd;
sos_loop[0].somModel.sram_ptr[6][577]=3;
sos_loop[0].somModel.sram_dat[6][578][0]=96'he4f1;
sos_loop[0].somModel.sram_ptr[6][578]=3;
sos_loop[0].somModel.sram_dat[6][579][0]=96'hd34e;
sos_loop[0].somModel.sram_ptr[6][579]=3;
sos_loop[0].somModel.sram_dat[6][580][0]=96'h28f9;
sos_loop[0].somModel.sram_ptr[6][580]=3;
sos_loop[0].somModel.sram_dat[6][581][0]=96'h7c60;
sos_loop[0].somModel.sram_ptr[6][581]=3;
sos_loop[0].somModel.sram_dat[6][582][0]=96'hd4d5;
sos_loop[0].somModel.sram_ptr[6][582]=3;
sos_loop[0].somModel.sram_dat[6][583][0]=96'h4278;
sos_loop[0].somModel.sram_ptr[6][583]=3;
sos_loop[0].somModel.sram_dat[6][584][0]=96'h2823;
sos_loop[0].somModel.sram_ptr[6][584]=3;
sos_loop[0].somModel.sram_dat[6][585][0]=96'hdf68;
sos_loop[0].somModel.sram_ptr[6][585]=3;
sos_loop[0].somModel.sram_dat[6][586][0]=96'h7947;
sos_loop[0].somModel.sram_ptr[6][586]=3;
sos_loop[0].somModel.sram_dat[6][587][0]=96'ha587;
sos_loop[0].somModel.sram_ptr[6][587]=3;
sos_loop[0].somModel.sram_dat[6][588][0]=96'h51ce;
sos_loop[0].somModel.sram_ptr[6][588]=3;
sos_loop[0].somModel.sram_dat[6][589][0]=96'h110a;
sos_loop[0].somModel.sram_ptr[6][589]=3;
sos_loop[0].somModel.sram_dat[6][590][0]=96'heffe;
sos_loop[0].somModel.sram_ptr[6][590]=3;
sos_loop[0].somModel.sram_dat[6][591][0]=96'hd97;
sos_loop[0].somModel.sram_ptr[6][591]=3;
sos_loop[0].somModel.sram_dat[6][592][0]=96'h2191;
sos_loop[0].somModel.sram_ptr[6][592]=3;
sos_loop[0].somModel.sram_dat[6][593][0]=96'ha878;
sos_loop[0].somModel.sram_ptr[6][593]=3;
sos_loop[0].somModel.sram_dat[6][594][0]=96'hf873;
sos_loop[0].somModel.sram_ptr[6][594]=3;
sos_loop[0].somModel.sram_dat[6][595][0]=96'hdf00;
sos_loop[0].somModel.sram_ptr[6][595]=3;
sos_loop[0].somModel.sram_dat[6][596][0]=96'h8139;
sos_loop[0].somModel.sram_ptr[6][596]=3;
sos_loop[0].somModel.sram_dat[6][597][0]=96'h5538;
sos_loop[0].somModel.sram_ptr[6][597]=3;
sos_loop[0].somModel.sram_dat[6][598][0]=96'he1ce;
sos_loop[0].somModel.sram_ptr[6][598]=3;
sos_loop[0].somModel.sram_dat[6][599][0]=96'h34dc;
sos_loop[0].somModel.sram_ptr[6][599]=3;
sos_loop[0].somModel.sram_dat[6][600][0]=96'h751e;
sos_loop[0].somModel.sram_ptr[6][600]=3;
sos_loop[0].somModel.sram_dat[6][601][0]=96'h48e3;
sos_loop[0].somModel.sram_ptr[6][601]=3;
sos_loop[0].somModel.sram_dat[6][602][0]=96'hd719;
sos_loop[0].somModel.sram_ptr[6][602]=3;
sos_loop[0].somModel.sram_dat[6][603][0]=96'h6f67;
sos_loop[0].somModel.sram_ptr[6][603]=3;
sos_loop[0].somModel.sram_dat[6][604][0]=96'hd5af;
sos_loop[0].somModel.sram_ptr[6][604]=3;
sos_loop[0].somModel.sram_dat[6][605][0]=96'h1c7c;
sos_loop[0].somModel.sram_ptr[6][605]=3;
sos_loop[0].somModel.sram_dat[6][606][0]=96'h5a36;
sos_loop[0].somModel.sram_ptr[6][606]=3;
sos_loop[0].somModel.sram_dat[6][607][0]=96'h5647;
sos_loop[0].somModel.sram_ptr[6][607]=3;
sos_loop[0].somModel.sram_dat[6][608][0]=96'ha79e;
sos_loop[0].somModel.sram_ptr[6][608]=3;
sos_loop[0].somModel.sram_dat[6][609][0]=96'hb278;
sos_loop[0].somModel.sram_ptr[6][609]=3;
sos_loop[0].somModel.sram_dat[6][610][0]=96'h40bf;
sos_loop[0].somModel.sram_ptr[6][610]=3;
sos_loop[0].somModel.sram_dat[6][611][0]=96'h799e;
sos_loop[0].somModel.sram_ptr[6][611]=3;
sos_loop[0].somModel.sram_dat[6][612][0]=96'hb51c;
sos_loop[0].somModel.sram_ptr[6][612]=3;
sos_loop[0].somModel.sram_dat[6][613][0]=96'heb9a;
sos_loop[0].somModel.sram_ptr[6][613]=3;
sos_loop[0].somModel.sram_dat[6][614][0]=96'h3e44;
sos_loop[0].somModel.sram_ptr[6][614]=3;
sos_loop[0].somModel.sram_dat[6][615][0]=96'h88bd;
sos_loop[0].somModel.sram_ptr[6][615]=3;
sos_loop[0].somModel.sram_dat[6][616][0]=96'h6126;
sos_loop[0].somModel.sram_ptr[6][616]=3;
sos_loop[0].somModel.sram_dat[6][617][0]=96'he67b;
sos_loop[0].somModel.sram_ptr[6][617]=3;
sos_loop[0].somModel.sram_dat[6][618][0]=96'hb998;
sos_loop[0].somModel.sram_ptr[6][618]=3;
sos_loop[0].somModel.sram_dat[6][619][0]=96'h82fe;
sos_loop[0].somModel.sram_ptr[6][619]=3;
sos_loop[0].somModel.sram_dat[6][620][0]=96'h3203;
sos_loop[0].somModel.sram_ptr[6][620]=3;
sos_loop[0].somModel.sram_dat[6][621][0]=96'hd92b;
sos_loop[0].somModel.sram_ptr[6][621]=3;
sos_loop[0].somModel.sram_dat[6][622][0]=96'h80ec;
sos_loop[0].somModel.sram_ptr[6][622]=3;
sos_loop[0].somModel.sram_dat[6][623][0]=96'h7aa1;
sos_loop[0].somModel.sram_ptr[6][623]=3;
sos_loop[0].somModel.sram_dat[6][624][0]=96'hfff3;
sos_loop[0].somModel.sram_ptr[6][624]=3;
sos_loop[0].somModel.sram_dat[6][625][0]=96'h19f1;
sos_loop[0].somModel.sram_ptr[6][625]=3;
sos_loop[0].somModel.sram_dat[6][626][0]=96'he2d3;
sos_loop[0].somModel.sram_ptr[6][626]=3;
sos_loop[0].somModel.sram_dat[6][627][0]=96'h1c4b;
sos_loop[0].somModel.sram_ptr[6][627]=3;
sos_loop[0].somModel.sram_dat[6][628][0]=96'hf785;
sos_loop[0].somModel.sram_ptr[6][628]=3;
sos_loop[0].somModel.sram_dat[6][629][0]=96'h6e92;
sos_loop[0].somModel.sram_ptr[6][629]=3;
sos_loop[0].somModel.sram_dat[6][630][0]=96'h8164;
sos_loop[0].somModel.sram_ptr[6][630]=3;
sos_loop[0].somModel.sram_dat[6][631][0]=96'hc136;
sos_loop[0].somModel.sram_ptr[6][631]=3;
sos_loop[0].somModel.sram_dat[6][632][0]=96'h79d2;
sos_loop[0].somModel.sram_ptr[6][632]=3;
sos_loop[0].somModel.sram_dat[6][633][0]=96'he175;
sos_loop[0].somModel.sram_ptr[6][633]=3;
sos_loop[0].somModel.sram_dat[6][634][0]=96'h6eda;
sos_loop[0].somModel.sram_ptr[6][634]=3;
sos_loop[0].somModel.sram_dat[6][635][0]=96'h6c68;
sos_loop[0].somModel.sram_ptr[6][635]=3;
sos_loop[0].somModel.sram_dat[6][636][0]=96'hbe89;
sos_loop[0].somModel.sram_ptr[6][636]=3;
sos_loop[0].somModel.sram_dat[6][637][0]=96'hd49f;
sos_loop[0].somModel.sram_ptr[6][637]=3;
sos_loop[0].somModel.sram_dat[6][638][0]=96'h9a7f;
sos_loop[0].somModel.sram_ptr[6][638]=3;
sos_loop[0].somModel.sram_dat[6][639][0]=96'h4960;
sos_loop[0].somModel.sram_ptr[6][639]=3;
sos_loop[0].somModel.sram_dat[6][640][0]=96'h1bc1;
sos_loop[0].somModel.sram_ptr[6][640]=3;
sos_loop[0].somModel.sram_dat[6][641][0]=96'h144e;
sos_loop[0].somModel.sram_ptr[6][641]=3;
sos_loop[0].somModel.sram_dat[6][642][0]=96'h779c;
sos_loop[0].somModel.sram_ptr[6][642]=3;
sos_loop[0].somModel.sram_dat[6][643][0]=96'h871a;
sos_loop[0].somModel.sram_ptr[6][643]=3;
sos_loop[0].somModel.sram_dat[6][644][0]=96'h1b85;
sos_loop[0].somModel.sram_ptr[6][644]=3;
sos_loop[0].somModel.sram_dat[6][645][0]=96'hb1e;
sos_loop[0].somModel.sram_ptr[6][645]=3;
sos_loop[0].somModel.sram_dat[6][646][0]=96'h573c;
sos_loop[0].somModel.sram_ptr[6][646]=3;
sos_loop[0].somModel.sram_dat[6][647][0]=96'h43ec;
sos_loop[0].somModel.sram_ptr[6][647]=3;
sos_loop[0].somModel.sram_dat[6][648][0]=96'h9e70;
sos_loop[0].somModel.sram_ptr[6][648]=3;
sos_loop[0].somModel.sram_dat[6][649][0]=96'h7bbb;
sos_loop[0].somModel.sram_ptr[6][649]=3;
sos_loop[0].somModel.sram_dat[6][650][0]=96'h58a8;
sos_loop[0].somModel.sram_ptr[6][650]=3;
sos_loop[0].somModel.sram_dat[6][651][0]=96'hbb95;
sos_loop[0].somModel.sram_ptr[6][651]=3;
sos_loop[0].somModel.sram_dat[6][652][0]=96'h4ee1;
sos_loop[0].somModel.sram_ptr[6][652]=3;
sos_loop[0].somModel.sram_dat[6][653][0]=96'hcd5e;
sos_loop[0].somModel.sram_ptr[6][653]=3;
sos_loop[0].somModel.sram_dat[6][654][0]=96'h855f;
sos_loop[0].somModel.sram_ptr[6][654]=3;
sos_loop[0].somModel.sram_dat[6][655][0]=96'h7a49;
sos_loop[0].somModel.sram_ptr[6][655]=3;
sos_loop[0].somModel.sram_dat[6][656][0]=96'h1c06;
sos_loop[0].somModel.sram_ptr[6][656]=3;
sos_loop[0].somModel.sram_dat[6][657][0]=96'hdc16;
sos_loop[0].somModel.sram_ptr[6][657]=3;
sos_loop[0].somModel.sram_dat[6][658][0]=96'h618d;
sos_loop[0].somModel.sram_ptr[6][658]=3;
sos_loop[0].somModel.sram_dat[6][659][0]=96'h7ea0;
sos_loop[0].somModel.sram_ptr[6][659]=3;
sos_loop[0].somModel.sram_dat[6][660][0]=96'hd910;
sos_loop[0].somModel.sram_ptr[6][660]=3;
sos_loop[0].somModel.sram_dat[6][661][0]=96'hdc31;
sos_loop[0].somModel.sram_ptr[6][661]=3;
sos_loop[0].somModel.sram_dat[6][662][0]=96'h88aa;
sos_loop[0].somModel.sram_ptr[6][662]=3;
sos_loop[0].somModel.sram_dat[6][663][0]=96'h89fe;
sos_loop[0].somModel.sram_ptr[6][663]=3;
sos_loop[0].somModel.sram_dat[6][664][0]=96'hf777;
sos_loop[0].somModel.sram_ptr[6][664]=3;
sos_loop[0].somModel.sram_dat[6][665][0]=96'h28d5;
sos_loop[0].somModel.sram_ptr[6][665]=3;
sos_loop[0].somModel.sram_dat[6][666][0]=96'h5497;
sos_loop[0].somModel.sram_ptr[6][666]=3;
sos_loop[0].somModel.sram_dat[6][667][0]=96'h9db1;
sos_loop[0].somModel.sram_ptr[6][667]=3;
sos_loop[0].somModel.sram_dat[6][668][0]=96'h570;
sos_loop[0].somModel.sram_ptr[6][668]=3;
sos_loop[0].somModel.sram_dat[6][669][0]=96'he79a;
sos_loop[0].somModel.sram_ptr[6][669]=3;
sos_loop[0].somModel.sram_dat[6][670][0]=96'haa71;
sos_loop[0].somModel.sram_ptr[6][670]=3;
sos_loop[0].somModel.sram_dat[6][671][0]=96'hdd36;
sos_loop[0].somModel.sram_ptr[6][671]=3;
sos_loop[0].somModel.sram_dat[6][672][0]=96'h77a3;
sos_loop[0].somModel.sram_ptr[6][672]=3;
sos_loop[0].somModel.sram_dat[6][673][0]=96'h2946;
sos_loop[0].somModel.sram_ptr[6][673]=3;
sos_loop[0].somModel.sram_dat[6][674][0]=96'hc3d1;
sos_loop[0].somModel.sram_ptr[6][674]=3;
sos_loop[0].somModel.sram_dat[6][675][0]=96'h884e;
sos_loop[0].somModel.sram_ptr[6][675]=3;
sos_loop[0].somModel.sram_dat[6][676][0]=96'h552c;
sos_loop[0].somModel.sram_ptr[6][676]=3;
sos_loop[0].somModel.sram_dat[6][677][0]=96'h418f;
sos_loop[0].somModel.sram_ptr[6][677]=3;
sos_loop[0].somModel.sram_dat[6][678][0]=96'h2d0;
sos_loop[0].somModel.sram_ptr[6][678]=3;
sos_loop[0].somModel.sram_dat[6][679][0]=96'h1688;
sos_loop[0].somModel.sram_ptr[6][679]=3;
sos_loop[0].somModel.sram_dat[6][680][0]=96'hd1ea;
sos_loop[0].somModel.sram_ptr[6][680]=3;
sos_loop[0].somModel.sram_dat[6][681][0]=96'hed72;
sos_loop[0].somModel.sram_ptr[6][681]=3;
sos_loop[0].somModel.sram_dat[6][682][0]=96'h4b54;
sos_loop[0].somModel.sram_ptr[6][682]=3;
sos_loop[0].somModel.sram_dat[6][683][0]=96'ha5ad;
sos_loop[0].somModel.sram_ptr[6][683]=3;
sos_loop[0].somModel.sram_dat[6][684][0]=96'h2270;
sos_loop[0].somModel.sram_ptr[6][684]=3;
sos_loop[0].somModel.sram_dat[6][685][0]=96'h7c75;
sos_loop[0].somModel.sram_ptr[6][685]=3;
sos_loop[0].somModel.sram_dat[6][686][0]=96'h3d8c;
sos_loop[0].somModel.sram_ptr[6][686]=3;
sos_loop[0].somModel.sram_dat[6][687][0]=96'h54cc;
sos_loop[0].somModel.sram_ptr[6][687]=3;
sos_loop[0].somModel.sram_dat[6][688][0]=96'h8f89;
sos_loop[0].somModel.sram_ptr[6][688]=3;
sos_loop[0].somModel.sram_dat[6][689][0]=96'h641e;
sos_loop[0].somModel.sram_ptr[6][689]=3;
sos_loop[0].somModel.sram_dat[6][690][0]=96'h66d;
sos_loop[0].somModel.sram_ptr[6][690]=3;
sos_loop[0].somModel.sram_dat[6][691][0]=96'hf56a;
sos_loop[0].somModel.sram_ptr[6][691]=3;
sos_loop[0].somModel.sram_dat[6][692][0]=96'h478;
sos_loop[0].somModel.sram_ptr[6][692]=3;
sos_loop[0].somModel.sram_dat[6][693][0]=96'h668d;
sos_loop[0].somModel.sram_ptr[6][693]=3;
sos_loop[0].somModel.sram_dat[6][694][0]=96'ha161;
sos_loop[0].somModel.sram_ptr[6][694]=3;
sos_loop[0].somModel.sram_dat[6][695][0]=96'h6b35;
sos_loop[0].somModel.sram_ptr[6][695]=3;
sos_loop[0].somModel.sram_dat[6][696][0]=96'h5b97;
sos_loop[0].somModel.sram_ptr[6][696]=3;
sos_loop[0].somModel.sram_dat[6][697][0]=96'hf63c;
sos_loop[0].somModel.sram_ptr[6][697]=3;
sos_loop[0].somModel.sram_dat[6][698][0]=96'h5629;
sos_loop[0].somModel.sram_ptr[6][698]=3;
sos_loop[0].somModel.sram_dat[6][699][0]=96'h2745;
sos_loop[0].somModel.sram_ptr[6][699]=3;
sos_loop[0].somModel.sram_dat[6][700][0]=96'h232e;
sos_loop[0].somModel.sram_ptr[6][700]=3;
sos_loop[0].somModel.cfg_tbl_sel[6] = 6;
sos_loop[0].somModel.cfg_dat_sel[6] = 0;
sos_loop[0].somModel.cfg_dat_vld[6] = 1;
sos_loop[0].somModel.cfg_miss_ptr[6] = 0;
sos_loop[0].somModel.tcam_data[7][0][0]=80'h00000000000000000000;
sos_loop[0].somModel.tcam_mask[7][0][0]=80'hffffffffffffffffffff;
sos_loop[0].somModel.tcam_data[7][1][0]=80'h00000000c76428a3ac18;
sos_loop[0].somModel.tcam_mask[7][1][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][2][0]=80'h000000006fa2b332a044;
sos_loop[0].somModel.tcam_mask[7][2][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][3][0]=80'h00000000df160ea7e244;
sos_loop[0].somModel.tcam_mask[7][3][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][4][0]=80'h00000000bde8a5158a2b;
sos_loop[0].somModel.tcam_mask[7][4][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][5][0]=80'h000000001c7fcaa5772f;
sos_loop[0].somModel.tcam_mask[7][5][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][6][0]=80'h00000000398bc2065413;
sos_loop[0].somModel.tcam_mask[7][6][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][7][0]=80'h00000000bf26a132d23e;
sos_loop[0].somModel.tcam_mask[7][7][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][8][0]=80'h000000002e5a52ddfb3f;
sos_loop[0].somModel.tcam_mask[7][8][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][9][0]=80'h000000000f9c4f448c4c;
sos_loop[0].somModel.tcam_mask[7][9][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][10][0]=80'h0000000035e4dd182f90;
sos_loop[0].somModel.tcam_mask[7][10][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][11][0]=80'h000000008513d0c50521;
sos_loop[0].somModel.tcam_mask[7][11][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][12][0]=80'h0000000035a66285b62e;
sos_loop[0].somModel.tcam_mask[7][12][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][13][0]=80'h000000004915d9de428f;
sos_loop[0].somModel.tcam_mask[7][13][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][14][0]=80'h000000003eff489073c2;
sos_loop[0].somModel.tcam_mask[7][14][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][15][0]=80'h00000000d00165db49c5;
sos_loop[0].somModel.tcam_mask[7][15][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][16][0]=80'h00000000c6e7d540048a;
sos_loop[0].somModel.tcam_mask[7][16][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][17][0]=80'h000000000d2cf31221e9;
sos_loop[0].somModel.tcam_mask[7][17][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][18][0]=80'h000000009cc2400c08bc;
sos_loop[0].somModel.tcam_mask[7][18][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][19][0]=80'h00000000e84ab68b1a24;
sos_loop[0].somModel.tcam_mask[7][19][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][20][0]=80'h00000000dc9c606e91ae;
sos_loop[0].somModel.tcam_mask[7][20][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][21][0]=80'h000000004b8ee53f7660;
sos_loop[0].somModel.tcam_mask[7][21][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][22][0]=80'h00000000a6dc109cdbbd;
sos_loop[0].somModel.tcam_mask[7][22][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][23][0]=80'h000000002e5acd726cb2;
sos_loop[0].somModel.tcam_mask[7][23][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][24][0]=80'h00000000bb30b2ecd487;
sos_loop[0].somModel.tcam_mask[7][24][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][25][0]=80'h000000009aeec82f8fac;
sos_loop[0].somModel.tcam_mask[7][25][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][26][0]=80'h00000000ab83fe2b985c;
sos_loop[0].somModel.tcam_mask[7][26][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][27][0]=80'h00000000ca3daac02b2f;
sos_loop[0].somModel.tcam_mask[7][27][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][28][0]=80'h000000001a893b2ffa10;
sos_loop[0].somModel.tcam_mask[7][28][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][29][0]=80'h00000000cb1ab883d9ca;
sos_loop[0].somModel.tcam_mask[7][29][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][30][0]=80'h000000006ddb0412e88d;
sos_loop[0].somModel.tcam_mask[7][30][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][31][0]=80'h0000000025d034a677c8;
sos_loop[0].somModel.tcam_mask[7][31][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][32][0]=80'h0000000002ee63ce89af;
sos_loop[0].somModel.tcam_mask[7][32][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[7][33][0]=80'h000000001ab5a710d843;
sos_loop[0].somModel.tcam_mask[7][33][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][34][0]=80'h0000000097e8c062f084;
sos_loop[0].somModel.tcam_mask[7][34][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][35][0]=80'h0000000030a809743d4f;
sos_loop[0].somModel.tcam_mask[7][35][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][36][0]=80'h0000000022420da7f8f4;
sos_loop[0].somModel.tcam_mask[7][36][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][37][0]=80'h00000000afaf284ad3bc;
sos_loop[0].somModel.tcam_mask[7][37][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][38][0]=80'h0000000053bd4f0d7794;
sos_loop[0].somModel.tcam_mask[7][38][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][39][0]=80'h000000005c0d39f2f061;
sos_loop[0].somModel.tcam_mask[7][39][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][40][0]=80'h000000009419a7ce074a;
sos_loop[0].somModel.tcam_mask[7][40][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][41][0]=80'h00000000052d45cc1e4a;
sos_loop[0].somModel.tcam_mask[7][41][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][42][0]=80'h000000009b30665b9971;
sos_loop[0].somModel.tcam_mask[7][42][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][43][0]=80'h0000000020d936f412c1;
sos_loop[0].somModel.tcam_mask[7][43][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][44][0]=80'h000000008b889af41550;
sos_loop[0].somModel.tcam_mask[7][44][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][45][0]=80'h00000000f91ce85e797d;
sos_loop[0].somModel.tcam_mask[7][45][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][46][0]=80'h0000000006e1dbd81191;
sos_loop[0].somModel.tcam_mask[7][46][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][47][0]=80'h00000000345e3c5f1365;
sos_loop[0].somModel.tcam_mask[7][47][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][48][0]=80'h000000008dceefe91dc9;
sos_loop[0].somModel.tcam_mask[7][48][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][49][0]=80'h00000000d47d2191ffed;
sos_loop[0].somModel.tcam_mask[7][49][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][50][0]=80'h000000007d341fbc821b;
sos_loop[0].somModel.tcam_mask[7][50][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][51][0]=80'h000000002e1c5d9ff7d9;
sos_loop[0].somModel.tcam_mask[7][51][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][52][0]=80'h00000000b7c667fd0324;
sos_loop[0].somModel.tcam_mask[7][52][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][53][0]=80'h000000004933bf21a16c;
sos_loop[0].somModel.tcam_mask[7][53][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][54][0]=80'h00000000f9724902347e;
sos_loop[0].somModel.tcam_mask[7][54][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][55][0]=80'h00000000aeb766b220db;
sos_loop[0].somModel.tcam_mask[7][55][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][56][0]=80'h00000000dbbc2a3224ab;
sos_loop[0].somModel.tcam_mask[7][56][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][57][0]=80'h00000000365a679e8085;
sos_loop[0].somModel.tcam_mask[7][57][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][58][0]=80'h00000000eeff7c2b7b33;
sos_loop[0].somModel.tcam_mask[7][58][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][59][0]=80'h0000000045bb6a31bb68;
sos_loop[0].somModel.tcam_mask[7][59][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][60][0]=80'h000000001a81b1c43f91;
sos_loop[0].somModel.tcam_mask[7][60][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][61][0]=80'h000000001de0ad29184a;
sos_loop[0].somModel.tcam_mask[7][61][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][62][0]=80'h000000004eb9229cd415;
sos_loop[0].somModel.tcam_mask[7][62][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][63][0]=80'h0000000075c39cfd15db;
sos_loop[0].somModel.tcam_mask[7][63][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][64][0]=80'h000000000bd7d9ddf726;
sos_loop[0].somModel.tcam_mask[7][64][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][65][0]=80'h00000000788ece7eed43;
sos_loop[0].somModel.tcam_mask[7][65][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][66][0]=80'h00000000689790000fff;
sos_loop[0].somModel.tcam_mask[7][66][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][67][0]=80'h0000000030fca31cf96b;
sos_loop[0].somModel.tcam_mask[7][67][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][68][0]=80'h00000000358975cc2823;
sos_loop[0].somModel.tcam_mask[7][68][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][69][0]=80'h000000006b1cd921c79d;
sos_loop[0].somModel.tcam_mask[7][69][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][70][0]=80'h00000000549a31ff63b7;
sos_loop[0].somModel.tcam_mask[7][70][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][71][0]=80'h00000000310dee607220;
sos_loop[0].somModel.tcam_mask[7][71][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][72][0]=80'h00000000af90fc2fb606;
sos_loop[0].somModel.tcam_mask[7][72][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][73][0]=80'h000000000db655000d3a;
sos_loop[0].somModel.tcam_mask[7][73][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][74][0]=80'h000000008bf35344ab45;
sos_loop[0].somModel.tcam_mask[7][74][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][75][0]=80'h000000002d8a38190b20;
sos_loop[0].somModel.tcam_mask[7][75][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][76][0]=80'h000000000263f7f66582;
sos_loop[0].somModel.tcam_mask[7][76][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[7][77][0]=80'h000000004dfc2ba4768d;
sos_loop[0].somModel.tcam_mask[7][77][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][78][0]=80'h00000000849983bfbe7a;
sos_loop[0].somModel.tcam_mask[7][78][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][79][0]=80'h000000001efcb2f4dd4d;
sos_loop[0].somModel.tcam_mask[7][79][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][80][0]=80'h0000000061e5a9de4569;
sos_loop[0].somModel.tcam_mask[7][80][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][81][0]=80'h00000000770c1c4bd3a5;
sos_loop[0].somModel.tcam_mask[7][81][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][82][0]=80'h00000000500562660aff;
sos_loop[0].somModel.tcam_mask[7][82][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][83][0]=80'h00000000a72a189143e2;
sos_loop[0].somModel.tcam_mask[7][83][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][84][0]=80'h0000000051a64abf0e09;
sos_loop[0].somModel.tcam_mask[7][84][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][85][0]=80'h000000001f5700abe928;
sos_loop[0].somModel.tcam_mask[7][85][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][86][0]=80'h00000000512e72fad6a2;
sos_loop[0].somModel.tcam_mask[7][86][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][87][0]=80'h000000005f3a530396cf;
sos_loop[0].somModel.tcam_mask[7][87][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][88][0]=80'h00000000748487400445;
sos_loop[0].somModel.tcam_mask[7][88][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][89][0]=80'h0000000087719fb3f864;
sos_loop[0].somModel.tcam_mask[7][89][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][90][0]=80'h00000000e88c8f60061d;
sos_loop[0].somModel.tcam_mask[7][90][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][91][0]=80'h000000009f6cc5f93019;
sos_loop[0].somModel.tcam_mask[7][91][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][92][0]=80'h00000000fa9df2c0fa11;
sos_loop[0].somModel.tcam_mask[7][92][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][93][0]=80'h000000003e5de237f4f3;
sos_loop[0].somModel.tcam_mask[7][93][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][94][0]=80'h000000001220e6f8b9fd;
sos_loop[0].somModel.tcam_mask[7][94][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][95][0]=80'h00000000ceb0c2f94c3c;
sos_loop[0].somModel.tcam_mask[7][95][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][96][0]=80'h000000001845b8356ded;
sos_loop[0].somModel.tcam_mask[7][96][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][97][0]=80'h00000000cb7d6f052ed9;
sos_loop[0].somModel.tcam_mask[7][97][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][98][0]=80'h00000000a1d827523dc7;
sos_loop[0].somModel.tcam_mask[7][98][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][99][0]=80'h000000000caf8264a3ea;
sos_loop[0].somModel.tcam_mask[7][99][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][100][0]=80'h0000000038ead3f12916;
sos_loop[0].somModel.tcam_mask[7][100][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][101][0]=80'h0000000013d2ee37c448;
sos_loop[0].somModel.tcam_mask[7][101][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][102][0]=80'h000000003c2fe7d9f34c;
sos_loop[0].somModel.tcam_mask[7][102][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][103][0]=80'h000000003c1db8626079;
sos_loop[0].somModel.tcam_mask[7][103][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][104][0]=80'h00000000865b861ca607;
sos_loop[0].somModel.tcam_mask[7][104][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][105][0]=80'h00000000794600c6d0f4;
sos_loop[0].somModel.tcam_mask[7][105][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][106][0]=80'h00000000e00c57f6e0b3;
sos_loop[0].somModel.tcam_mask[7][106][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][107][0]=80'h00000000e29db65e8903;
sos_loop[0].somModel.tcam_mask[7][107][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][108][0]=80'h000000008e261e6170f3;
sos_loop[0].somModel.tcam_mask[7][108][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][109][0]=80'h0000000066939b10ec73;
sos_loop[0].somModel.tcam_mask[7][109][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][110][0]=80'h0000000070c2e9c3c8eb;
sos_loop[0].somModel.tcam_mask[7][110][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][111][0]=80'h0000000045c66be84cf4;
sos_loop[0].somModel.tcam_mask[7][111][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][112][0]=80'h00000000232cef211d0e;
sos_loop[0].somModel.tcam_mask[7][112][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][113][0]=80'h0000000080542dda5aa2;
sos_loop[0].somModel.tcam_mask[7][113][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][114][0]=80'h00000000474effbc30dd;
sos_loop[0].somModel.tcam_mask[7][114][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][115][0]=80'h00000000e4cebd5c6fa4;
sos_loop[0].somModel.tcam_mask[7][115][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][116][0]=80'h00000000af6a54830375;
sos_loop[0].somModel.tcam_mask[7][116][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][117][0]=80'h000000008ef028be44c1;
sos_loop[0].somModel.tcam_mask[7][117][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][118][0]=80'h000000005fdca8436bf4;
sos_loop[0].somModel.tcam_mask[7][118][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][119][0]=80'h000000006e7e1c15bd08;
sos_loop[0].somModel.tcam_mask[7][119][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][120][0]=80'h00000000134c1f65fd66;
sos_loop[0].somModel.tcam_mask[7][120][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][121][0]=80'h00000000cea87493679f;
sos_loop[0].somModel.tcam_mask[7][121][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][122][0]=80'h00000000ceb7bc309c1a;
sos_loop[0].somModel.tcam_mask[7][122][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][123][0]=80'h0000000061a6f8771878;
sos_loop[0].somModel.tcam_mask[7][123][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][124][0]=80'h00000000cedef6a567fe;
sos_loop[0].somModel.tcam_mask[7][124][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][125][0]=80'h000000002e32a08622cd;
sos_loop[0].somModel.tcam_mask[7][125][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][126][0]=80'h000000005356e16b8fd7;
sos_loop[0].somModel.tcam_mask[7][126][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][127][0]=80'h00000000fd605bd942c3;
sos_loop[0].somModel.tcam_mask[7][127][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][128][0]=80'h0000000000d5f103f449;
sos_loop[0].somModel.tcam_mask[7][128][0]=80'hffffffffff0000000000;
sos_loop[0].somModel.tcam_data[7][129][0]=80'h000000005f57f4362b22;
sos_loop[0].somModel.tcam_mask[7][129][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][130][0]=80'h000000002e67f284f871;
sos_loop[0].somModel.tcam_mask[7][130][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][131][0]=80'h00000000ecd79dcadc01;
sos_loop[0].somModel.tcam_mask[7][131][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][132][0]=80'h00000000e00525c7b0f8;
sos_loop[0].somModel.tcam_mask[7][132][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][133][0]=80'h00000000b3cf483e6c80;
sos_loop[0].somModel.tcam_mask[7][133][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][134][0]=80'h0000000077eb26f31bbe;
sos_loop[0].somModel.tcam_mask[7][134][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][135][0]=80'h000000008b676c49d915;
sos_loop[0].somModel.tcam_mask[7][135][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][136][0]=80'h000000000a2822acbd35;
sos_loop[0].somModel.tcam_mask[7][136][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][137][0]=80'h0000000003a257929df1;
sos_loop[0].somModel.tcam_mask[7][137][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[7][138][0]=80'h00000000e9b0e1c40a18;
sos_loop[0].somModel.tcam_mask[7][138][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][139][0]=80'h000000003f10a0b32f42;
sos_loop[0].somModel.tcam_mask[7][139][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][140][0]=80'h00000000f8a042a8b1d1;
sos_loop[0].somModel.tcam_mask[7][140][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][141][0]=80'h00000000c010041f98fe;
sos_loop[0].somModel.tcam_mask[7][141][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][142][0]=80'h000000006f5155d6bf2a;
sos_loop[0].somModel.tcam_mask[7][142][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][143][0]=80'h000000006174e0aee88e;
sos_loop[0].somModel.tcam_mask[7][143][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][144][0]=80'h00000000d8f296505931;
sos_loop[0].somModel.tcam_mask[7][144][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][145][0]=80'h00000000e512e3c64789;
sos_loop[0].somModel.tcam_mask[7][145][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][146][0]=80'h00000000373e0b9976b9;
sos_loop[0].somModel.tcam_mask[7][146][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][147][0]=80'h0000000003e7dacda18b;
sos_loop[0].somModel.tcam_mask[7][147][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[7][148][0]=80'h000000000964ddbc00a5;
sos_loop[0].somModel.tcam_mask[7][148][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][149][0]=80'h0000000054781b947c65;
sos_loop[0].somModel.tcam_mask[7][149][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][150][0]=80'h000000004e476ae23070;
sos_loop[0].somModel.tcam_mask[7][150][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][151][0]=80'h00000000965a202c5dd1;
sos_loop[0].somModel.tcam_mask[7][151][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][152][0]=80'h000000006eeef25e5a0e;
sos_loop[0].somModel.tcam_mask[7][152][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][153][0]=80'h00000000bd9be825e53c;
sos_loop[0].somModel.tcam_mask[7][153][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][154][0]=80'h000000005a0d2b0e2652;
sos_loop[0].somModel.tcam_mask[7][154][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][155][0]=80'h00000000f02c2960a78f;
sos_loop[0].somModel.tcam_mask[7][155][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][156][0]=80'h0000000043801573ed5c;
sos_loop[0].somModel.tcam_mask[7][156][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][157][0]=80'h0000000034d1a3628645;
sos_loop[0].somModel.tcam_mask[7][157][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][158][0]=80'h00000000476d2c7ebc16;
sos_loop[0].somModel.tcam_mask[7][158][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][159][0]=80'h00000000a17de6c9b9c6;
sos_loop[0].somModel.tcam_mask[7][159][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][160][0]=80'h000000002e3b2da7cb0e;
sos_loop[0].somModel.tcam_mask[7][160][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][161][0]=80'h00000000618fe75b3a00;
sos_loop[0].somModel.tcam_mask[7][161][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][162][0]=80'h000000007868e9b929a2;
sos_loop[0].somModel.tcam_mask[7][162][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][163][0]=80'h00000000cbe5e4137d1a;
sos_loop[0].somModel.tcam_mask[7][163][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][164][0]=80'h000000006771e8c490b5;
sos_loop[0].somModel.tcam_mask[7][164][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][165][0]=80'h000000007be9cc15dbad;
sos_loop[0].somModel.tcam_mask[7][165][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][166][0]=80'h000000008c89b097b14c;
sos_loop[0].somModel.tcam_mask[7][166][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][167][0]=80'h00000000f2124342ae18;
sos_loop[0].somModel.tcam_mask[7][167][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][168][0]=80'h00000000330261ba3670;
sos_loop[0].somModel.tcam_mask[7][168][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][169][0]=80'h0000000042c4edb6d896;
sos_loop[0].somModel.tcam_mask[7][169][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][170][0]=80'h0000000023a570bc32da;
sos_loop[0].somModel.tcam_mask[7][170][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][171][0]=80'h00000000db4f2973fc73;
sos_loop[0].somModel.tcam_mask[7][171][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][172][0]=80'h000000004c40d88318b1;
sos_loop[0].somModel.tcam_mask[7][172][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][173][0]=80'h000000001273739101e3;
sos_loop[0].somModel.tcam_mask[7][173][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][174][0]=80'h000000009c2ebac8770d;
sos_loop[0].somModel.tcam_mask[7][174][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][175][0]=80'h00000000aaeaffde1744;
sos_loop[0].somModel.tcam_mask[7][175][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][176][0]=80'h0000000067b1d0406ac4;
sos_loop[0].somModel.tcam_mask[7][176][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][177][0]=80'h00000000602be7c25423;
sos_loop[0].somModel.tcam_mask[7][177][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][178][0]=80'h000000007bd2374d89da;
sos_loop[0].somModel.tcam_mask[7][178][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][179][0]=80'h00000000484efbf68ee5;
sos_loop[0].somModel.tcam_mask[7][179][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][180][0]=80'h000000008c2970d5df55;
sos_loop[0].somModel.tcam_mask[7][180][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][181][0]=80'h00000000aec65cebfe7b;
sos_loop[0].somModel.tcam_mask[7][181][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][182][0]=80'h0000000094dfc4cad63a;
sos_loop[0].somModel.tcam_mask[7][182][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][183][0]=80'h0000000016398c9c5329;
sos_loop[0].somModel.tcam_mask[7][183][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][184][0]=80'h00000000c1d9c5b84501;
sos_loop[0].somModel.tcam_mask[7][184][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][185][0]=80'h00000000d1ad3332662b;
sos_loop[0].somModel.tcam_mask[7][185][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][186][0]=80'h00000000b91d094ca5fa;
sos_loop[0].somModel.tcam_mask[7][186][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][187][0]=80'h0000000066807169ce5b;
sos_loop[0].somModel.tcam_mask[7][187][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][188][0]=80'h000000006ef096e4f564;
sos_loop[0].somModel.tcam_mask[7][188][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][189][0]=80'h00000000328864e675f7;
sos_loop[0].somModel.tcam_mask[7][189][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][190][0]=80'h000000007dae2b0e1b45;
sos_loop[0].somModel.tcam_mask[7][190][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][191][0]=80'h00000000bcb94b47b6e1;
sos_loop[0].somModel.tcam_mask[7][191][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][192][0]=80'h00000000969630df4be5;
sos_loop[0].somModel.tcam_mask[7][192][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][193][0]=80'h000000008fa1021a531a;
sos_loop[0].somModel.tcam_mask[7][193][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][194][0]=80'h00000000872d61d5debf;
sos_loop[0].somModel.tcam_mask[7][194][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][195][0]=80'h00000000991610788933;
sos_loop[0].somModel.tcam_mask[7][195][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][196][0]=80'h000000000abf899e0a35;
sos_loop[0].somModel.tcam_mask[7][196][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][197][0]=80'h000000009a50b37b4c4e;
sos_loop[0].somModel.tcam_mask[7][197][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][198][0]=80'h00000000a57859f9c477;
sos_loop[0].somModel.tcam_mask[7][198][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][199][0]=80'h000000000079cd60c49c;
sos_loop[0].somModel.tcam_mask[7][199][0]=80'hffffffffff8000000000;
sos_loop[0].somModel.tcam_data[7][200][0]=80'h00000000116a5a1abd7d;
sos_loop[0].somModel.tcam_mask[7][200][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][201][0]=80'h00000000c21fd0b46818;
sos_loop[0].somModel.tcam_mask[7][201][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][202][0]=80'h00000000cb7c1d8cfffa;
sos_loop[0].somModel.tcam_mask[7][202][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][203][0]=80'h000000005da2668e789f;
sos_loop[0].somModel.tcam_mask[7][203][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][204][0]=80'h00000000a975554d1660;
sos_loop[0].somModel.tcam_mask[7][204][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][205][0]=80'h00000000f527f8412a24;
sos_loop[0].somModel.tcam_mask[7][205][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][206][0]=80'h000000006e7cabe12a47;
sos_loop[0].somModel.tcam_mask[7][206][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][207][0]=80'h00000000ecce1c4cd86e;
sos_loop[0].somModel.tcam_mask[7][207][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][208][0]=80'h0000000072d3d3fcd72b;
sos_loop[0].somModel.tcam_mask[7][208][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][209][0]=80'h00000000839e1fb55d44;
sos_loop[0].somModel.tcam_mask[7][209][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][210][0]=80'h00000000478398e0b9ee;
sos_loop[0].somModel.tcam_mask[7][210][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][211][0]=80'h000000008530d50e759f;
sos_loop[0].somModel.tcam_mask[7][211][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][212][0]=80'h0000000011f968361ebd;
sos_loop[0].somModel.tcam_mask[7][212][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][213][0]=80'h000000008ce994cc083f;
sos_loop[0].somModel.tcam_mask[7][213][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][214][0]=80'h000000002c23f84988ee;
sos_loop[0].somModel.tcam_mask[7][214][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][215][0]=80'h000000009760938f25c2;
sos_loop[0].somModel.tcam_mask[7][215][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][216][0]=80'h00000000274efbfa8211;
sos_loop[0].somModel.tcam_mask[7][216][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][217][0]=80'h00000000694132b93ba3;
sos_loop[0].somModel.tcam_mask[7][217][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][218][0]=80'h000000000682f3056401;
sos_loop[0].somModel.tcam_mask[7][218][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][219][0]=80'h00000000d1c36a785d4f;
sos_loop[0].somModel.tcam_mask[7][219][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][220][0]=80'h000000004ae9b6d2ef4f;
sos_loop[0].somModel.tcam_mask[7][220][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][221][0]=80'h00000000c9c32ab41eeb;
sos_loop[0].somModel.tcam_mask[7][221][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][222][0]=80'h00000000cbc076ebe28e;
sos_loop[0].somModel.tcam_mask[7][222][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][223][0]=80'h00000000fbda31fd76c0;
sos_loop[0].somModel.tcam_mask[7][223][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][224][0]=80'h000000009a099a151b35;
sos_loop[0].somModel.tcam_mask[7][224][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][225][0]=80'h0000000054a1681b3ffb;
sos_loop[0].somModel.tcam_mask[7][225][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][226][0]=80'h00000000f0cf8f9ee272;
sos_loop[0].somModel.tcam_mask[7][226][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][227][0]=80'h000000003f535b44d28a;
sos_loop[0].somModel.tcam_mask[7][227][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][228][0]=80'h000000007ae44fa333c8;
sos_loop[0].somModel.tcam_mask[7][228][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][229][0]=80'h00000000b665ce7f735a;
sos_loop[0].somModel.tcam_mask[7][229][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][230][0]=80'h00000000626c7ae8774d;
sos_loop[0].somModel.tcam_mask[7][230][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][231][0]=80'h00000000f3cddb51d392;
sos_loop[0].somModel.tcam_mask[7][231][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][232][0]=80'h00000000944a75a8319c;
sos_loop[0].somModel.tcam_mask[7][232][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][233][0]=80'h00000000eaacb9890fae;
sos_loop[0].somModel.tcam_mask[7][233][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][234][0]=80'h00000000046f6540ec7f;
sos_loop[0].somModel.tcam_mask[7][234][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][235][0]=80'h00000000c6088fc1bd3d;
sos_loop[0].somModel.tcam_mask[7][235][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][236][0]=80'h000000005e0b61c56031;
sos_loop[0].somModel.tcam_mask[7][236][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][237][0]=80'h00000000027b4c51c3bb;
sos_loop[0].somModel.tcam_mask[7][237][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[7][238][0]=80'h00000000be4d82d7e60e;
sos_loop[0].somModel.tcam_mask[7][238][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][239][0]=80'h000000007eef6a0932c5;
sos_loop[0].somModel.tcam_mask[7][239][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][240][0]=80'h00000000564f40cb3bc6;
sos_loop[0].somModel.tcam_mask[7][240][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][241][0]=80'h0000000049ba0e14ede1;
sos_loop[0].somModel.tcam_mask[7][241][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][242][0]=80'h000000000ffa1385e8e1;
sos_loop[0].somModel.tcam_mask[7][242][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][243][0]=80'h00000000c2a6a6c5875c;
sos_loop[0].somModel.tcam_mask[7][243][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][244][0]=80'h0000000046ed88992ff9;
sos_loop[0].somModel.tcam_mask[7][244][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][245][0]=80'h000000007bd52c488741;
sos_loop[0].somModel.tcam_mask[7][245][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][246][0]=80'h00000000dd037b320186;
sos_loop[0].somModel.tcam_mask[7][246][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][247][0]=80'h00000000bc45bae8ac0a;
sos_loop[0].somModel.tcam_mask[7][247][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][248][0]=80'h000000005b06c7e96f30;
sos_loop[0].somModel.tcam_mask[7][248][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][249][0]=80'h00000000d4ddc557a673;
sos_loop[0].somModel.tcam_mask[7][249][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][250][0]=80'h0000000053ec21af6aa7;
sos_loop[0].somModel.tcam_mask[7][250][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][251][0]=80'h0000000017ac57f88e87;
sos_loop[0].somModel.tcam_mask[7][251][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][252][0]=80'h00000000a4100e4032cc;
sos_loop[0].somModel.tcam_mask[7][252][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][253][0]=80'h00000000140fa51dda60;
sos_loop[0].somModel.tcam_mask[7][253][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][254][0]=80'h00000000ba76b63b04af;
sos_loop[0].somModel.tcam_mask[7][254][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][255][0]=80'h000000007bf30212d42d;
sos_loop[0].somModel.tcam_mask[7][255][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][256][0]=80'h00000000389a856d0929;
sos_loop[0].somModel.tcam_mask[7][256][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][257][0]=80'h00000000971def77bfa0;
sos_loop[0].somModel.tcam_mask[7][257][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][258][0]=80'h000000007fea6ca2dda9;
sos_loop[0].somModel.tcam_mask[7][258][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][259][0]=80'h000000006cc87b7163e1;
sos_loop[0].somModel.tcam_mask[7][259][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][260][0]=80'h00000000652f37432033;
sos_loop[0].somModel.tcam_mask[7][260][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][261][0]=80'h0000000094ca0afeaf40;
sos_loop[0].somModel.tcam_mask[7][261][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][262][0]=80'h00000000aa6075a82cfd;
sos_loop[0].somModel.tcam_mask[7][262][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][263][0]=80'h00000000e393132fbd4d;
sos_loop[0].somModel.tcam_mask[7][263][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][264][0]=80'h000000008617fb8769a3;
sos_loop[0].somModel.tcam_mask[7][264][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][265][0]=80'h00000000d45704f554fa;
sos_loop[0].somModel.tcam_mask[7][265][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][266][0]=80'h00000000083aeac67707;
sos_loop[0].somModel.tcam_mask[7][266][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][267][0]=80'h00000000ad11dd592c9a;
sos_loop[0].somModel.tcam_mask[7][267][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][268][0]=80'h00000000199fcd09ed28;
sos_loop[0].somModel.tcam_mask[7][268][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][269][0]=80'h00000000306fc67d4fd2;
sos_loop[0].somModel.tcam_mask[7][269][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][270][0]=80'h00000000ded308236673;
sos_loop[0].somModel.tcam_mask[7][270][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][271][0]=80'h000000006bb4f3981543;
sos_loop[0].somModel.tcam_mask[7][271][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][272][0]=80'h0000000028d774fa8bab;
sos_loop[0].somModel.tcam_mask[7][272][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][273][0]=80'h000000005f39e126fa40;
sos_loop[0].somModel.tcam_mask[7][273][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][274][0]=80'h000000004ec1930dd830;
sos_loop[0].somModel.tcam_mask[7][274][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][275][0]=80'h000000002eabafa47444;
sos_loop[0].somModel.tcam_mask[7][275][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][276][0]=80'h00000000f2c4354979b5;
sos_loop[0].somModel.tcam_mask[7][276][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][277][0]=80'h000000004375ff2839ff;
sos_loop[0].somModel.tcam_mask[7][277][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][278][0]=80'h00000000831847d750e3;
sos_loop[0].somModel.tcam_mask[7][278][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][279][0]=80'h000000006d4ff70a7fc3;
sos_loop[0].somModel.tcam_mask[7][279][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][280][0]=80'h0000000067633ad96690;
sos_loop[0].somModel.tcam_mask[7][280][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][281][0]=80'h0000000058b1bb7ab35b;
sos_loop[0].somModel.tcam_mask[7][281][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][282][0]=80'h00000000378d65b1297a;
sos_loop[0].somModel.tcam_mask[7][282][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][283][0]=80'h000000008ab24a720a34;
sos_loop[0].somModel.tcam_mask[7][283][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][284][0]=80'h000000009b617faf808a;
sos_loop[0].somModel.tcam_mask[7][284][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][285][0]=80'h000000002b5be33345f9;
sos_loop[0].somModel.tcam_mask[7][285][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][286][0]=80'h0000000080b069925240;
sos_loop[0].somModel.tcam_mask[7][286][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][287][0]=80'h0000000064819ae5ce38;
sos_loop[0].somModel.tcam_mask[7][287][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][288][0]=80'h00000000c8a2886319ad;
sos_loop[0].somModel.tcam_mask[7][288][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][289][0]=80'h00000000bba80680cd74;
sos_loop[0].somModel.tcam_mask[7][289][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][290][0]=80'h00000000c624c1780420;
sos_loop[0].somModel.tcam_mask[7][290][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][291][0]=80'h000000000df4dc19f8a0;
sos_loop[0].somModel.tcam_mask[7][291][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][292][0]=80'h00000000bf4fc4c5109d;
sos_loop[0].somModel.tcam_mask[7][292][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][293][0]=80'h00000000230e53a6e40d;
sos_loop[0].somModel.tcam_mask[7][293][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][294][0]=80'h000000006a8845704812;
sos_loop[0].somModel.tcam_mask[7][294][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][295][0]=80'h00000000d02d7e61c3ff;
sos_loop[0].somModel.tcam_mask[7][295][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][296][0]=80'h0000000042d9ad4b7cb5;
sos_loop[0].somModel.tcam_mask[7][296][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][297][0]=80'h000000006620c43e40cd;
sos_loop[0].somModel.tcam_mask[7][297][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][298][0]=80'h00000000572b2a5075a9;
sos_loop[0].somModel.tcam_mask[7][298][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][299][0]=80'h000000000bc0a3cd8632;
sos_loop[0].somModel.tcam_mask[7][299][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][300][0]=80'h00000000318840f45c23;
sos_loop[0].somModel.tcam_mask[7][300][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][301][0]=80'h000000007ec0b9f2df84;
sos_loop[0].somModel.tcam_mask[7][301][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][302][0]=80'h000000000708eaeea371;
sos_loop[0].somModel.tcam_mask[7][302][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][303][0]=80'h0000000029e3e9901c1f;
sos_loop[0].somModel.tcam_mask[7][303][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][304][0]=80'h00000000f4f0fb40376f;
sos_loop[0].somModel.tcam_mask[7][304][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][305][0]=80'h000000007de8c27c7bf8;
sos_loop[0].somModel.tcam_mask[7][305][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][306][0]=80'h00000000722214538bb3;
sos_loop[0].somModel.tcam_mask[7][306][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][307][0]=80'h00000000b35284a2e8f3;
sos_loop[0].somModel.tcam_mask[7][307][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][308][0]=80'h00000000c1e963dc4088;
sos_loop[0].somModel.tcam_mask[7][308][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][309][0]=80'h0000000050d5503770e6;
sos_loop[0].somModel.tcam_mask[7][309][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][310][0]=80'h00000000b63951662a30;
sos_loop[0].somModel.tcam_mask[7][310][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][311][0]=80'h000000007eddea567619;
sos_loop[0].somModel.tcam_mask[7][311][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][312][0]=80'h000000004eab0a109e8f;
sos_loop[0].somModel.tcam_mask[7][312][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][313][0]=80'h00000000e549f26a551a;
sos_loop[0].somModel.tcam_mask[7][313][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][314][0]=80'h00000000161e12d7d5f4;
sos_loop[0].somModel.tcam_mask[7][314][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][315][0]=80'h000000002fb8691cf03d;
sos_loop[0].somModel.tcam_mask[7][315][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][316][0]=80'h000000006d0dd414bd88;
sos_loop[0].somModel.tcam_mask[7][316][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][317][0]=80'h00000000d47f0cfd8269;
sos_loop[0].somModel.tcam_mask[7][317][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][318][0]=80'h00000000e7fe58f76aac;
sos_loop[0].somModel.tcam_mask[7][318][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][319][0]=80'h00000000cddb5437e4b9;
sos_loop[0].somModel.tcam_mask[7][319][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][320][0]=80'h0000000058ac2d7d65c1;
sos_loop[0].somModel.tcam_mask[7][320][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][321][0]=80'h00000000e81d8eb85034;
sos_loop[0].somModel.tcam_mask[7][321][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][322][0]=80'h00000000a6fb99d69d1b;
sos_loop[0].somModel.tcam_mask[7][322][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][323][0]=80'h0000000085db0f2ad52e;
sos_loop[0].somModel.tcam_mask[7][323][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][324][0]=80'h00000000ba447f49c0b1;
sos_loop[0].somModel.tcam_mask[7][324][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][325][0]=80'h0000000099d3496acd35;
sos_loop[0].somModel.tcam_mask[7][325][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][326][0]=80'h0000000040e7e1b07303;
sos_loop[0].somModel.tcam_mask[7][326][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][327][0]=80'h0000000055f948ebe91d;
sos_loop[0].somModel.tcam_mask[7][327][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][328][0]=80'h00000000392c0459ce02;
sos_loop[0].somModel.tcam_mask[7][328][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][329][0]=80'h000000007e3d419f5d34;
sos_loop[0].somModel.tcam_mask[7][329][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][330][0]=80'h00000000e74efb58eaa7;
sos_loop[0].somModel.tcam_mask[7][330][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][331][0]=80'h00000000f83f581e4482;
sos_loop[0].somModel.tcam_mask[7][331][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][332][0]=80'h000000009cce1dfeef14;
sos_loop[0].somModel.tcam_mask[7][332][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][333][0]=80'h000000004b70936e9f64;
sos_loop[0].somModel.tcam_mask[7][333][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][334][0]=80'h000000008f60bf446783;
sos_loop[0].somModel.tcam_mask[7][334][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][335][0]=80'h0000000093a9046448e2;
sos_loop[0].somModel.tcam_mask[7][335][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][336][0]=80'h000000006e3ce4ac6730;
sos_loop[0].somModel.tcam_mask[7][336][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][337][0]=80'h0000000084de22fbc40a;
sos_loop[0].somModel.tcam_mask[7][337][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][338][0]=80'h000000002d98732c0914;
sos_loop[0].somModel.tcam_mask[7][338][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][339][0]=80'h00000000588e0584287c;
sos_loop[0].somModel.tcam_mask[7][339][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][340][0]=80'h000000008f50e0497e89;
sos_loop[0].somModel.tcam_mask[7][340][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][341][0]=80'h00000000b0e119fb2555;
sos_loop[0].somModel.tcam_mask[7][341][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][342][0]=80'h000000004cd3c2cde21a;
sos_loop[0].somModel.tcam_mask[7][342][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][343][0]=80'h00000000da342cb3beee;
sos_loop[0].somModel.tcam_mask[7][343][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][344][0]=80'h000000009f7fc5e6a042;
sos_loop[0].somModel.tcam_mask[7][344][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][345][0]=80'h00000000cc5300c82669;
sos_loop[0].somModel.tcam_mask[7][345][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][346][0]=80'h000000006a1ec386bf00;
sos_loop[0].somModel.tcam_mask[7][346][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][347][0]=80'h000000002317e8d90545;
sos_loop[0].somModel.tcam_mask[7][347][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][348][0]=80'h000000008d4fe98625cf;
sos_loop[0].somModel.tcam_mask[7][348][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][349][0]=80'h00000000060665e2c19e;
sos_loop[0].somModel.tcam_mask[7][349][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][350][0]=80'h00000000596674fbbfb1;
sos_loop[0].somModel.tcam_mask[7][350][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][351][0]=80'h000000005c7688d8aad5;
sos_loop[0].somModel.tcam_mask[7][351][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][352][0]=80'h0000000099c3cb202d30;
sos_loop[0].somModel.tcam_mask[7][352][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][353][0]=80'h00000000a86ac83a7681;
sos_loop[0].somModel.tcam_mask[7][353][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][354][0]=80'h00000000f9f330aaf7e5;
sos_loop[0].somModel.tcam_mask[7][354][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][355][0]=80'h000000003c3dcdb988e5;
sos_loop[0].somModel.tcam_mask[7][355][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][356][0]=80'h0000000082440e73e0a4;
sos_loop[0].somModel.tcam_mask[7][356][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][357][0]=80'h00000000deb63d376bdd;
sos_loop[0].somModel.tcam_mask[7][357][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][358][0]=80'h000000003f13c6d986da;
sos_loop[0].somModel.tcam_mask[7][358][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][359][0]=80'h00000000959a11161a8a;
sos_loop[0].somModel.tcam_mask[7][359][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][360][0]=80'h0000000004fc4b9709a2;
sos_loop[0].somModel.tcam_mask[7][360][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][361][0]=80'h000000000603260a4fa8;
sos_loop[0].somModel.tcam_mask[7][361][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][362][0]=80'h00000000317642426d30;
sos_loop[0].somModel.tcam_mask[7][362][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][363][0]=80'h0000000093eea5159da0;
sos_loop[0].somModel.tcam_mask[7][363][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][364][0]=80'h00000000a6a6c5effbb8;
sos_loop[0].somModel.tcam_mask[7][364][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][365][0]=80'h000000009a556fc0f1e1;
sos_loop[0].somModel.tcam_mask[7][365][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][366][0]=80'h00000000ca8bfde422b1;
sos_loop[0].somModel.tcam_mask[7][366][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][367][0]=80'h000000006b3d4da4a0e4;
sos_loop[0].somModel.tcam_mask[7][367][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][368][0]=80'h00000000b8725432eee0;
sos_loop[0].somModel.tcam_mask[7][368][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][369][0]=80'h000000002a5f4d97572c;
sos_loop[0].somModel.tcam_mask[7][369][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][370][0]=80'h0000000003f4b2f37c91;
sos_loop[0].somModel.tcam_mask[7][370][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[7][371][0]=80'h000000006d012a56f306;
sos_loop[0].somModel.tcam_mask[7][371][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][372][0]=80'h00000000f39c18ff7423;
sos_loop[0].somModel.tcam_mask[7][372][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][373][0]=80'h0000000064fe54c3d020;
sos_loop[0].somModel.tcam_mask[7][373][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][374][0]=80'h000000005941386df853;
sos_loop[0].somModel.tcam_mask[7][374][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][375][0]=80'h00000000fd5081a7023d;
sos_loop[0].somModel.tcam_mask[7][375][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][376][0]=80'h0000000059d252677e44;
sos_loop[0].somModel.tcam_mask[7][376][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][377][0]=80'h00000000b1ef710456c8;
sos_loop[0].somModel.tcam_mask[7][377][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][378][0]=80'h000000008a3b29afa55f;
sos_loop[0].somModel.tcam_mask[7][378][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][379][0]=80'h00000000a8f4af7c920a;
sos_loop[0].somModel.tcam_mask[7][379][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][380][0]=80'h000000009b5b556528f0;
sos_loop[0].somModel.tcam_mask[7][380][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][381][0]=80'h000000008d75c4ce6384;
sos_loop[0].somModel.tcam_mask[7][381][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][382][0]=80'h00000000644e172a4d39;
sos_loop[0].somModel.tcam_mask[7][382][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][383][0]=80'h000000004e2c31c4e9bf;
sos_loop[0].somModel.tcam_mask[7][383][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][384][0]=80'h00000000fb16e104670e;
sos_loop[0].somModel.tcam_mask[7][384][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][385][0]=80'h00000000edda66338267;
sos_loop[0].somModel.tcam_mask[7][385][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][386][0]=80'h00000000028c12a16f1b;
sos_loop[0].somModel.tcam_mask[7][386][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[7][387][0]=80'h00000000ff84824ad314;
sos_loop[0].somModel.tcam_mask[7][387][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][388][0]=80'h000000000be7756aeeab;
sos_loop[0].somModel.tcam_mask[7][388][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][389][0]=80'h000000007e61e055303f;
sos_loop[0].somModel.tcam_mask[7][389][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][390][0]=80'h00000000aac7193a22af;
sos_loop[0].somModel.tcam_mask[7][390][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][391][0]=80'h00000000565f0106873e;
sos_loop[0].somModel.tcam_mask[7][391][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][392][0]=80'h0000000075032e61802d;
sos_loop[0].somModel.tcam_mask[7][392][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][393][0]=80'h00000000f2f7c9dbbf6e;
sos_loop[0].somModel.tcam_mask[7][393][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][394][0]=80'h00000000c616b82074dc;
sos_loop[0].somModel.tcam_mask[7][394][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][395][0]=80'h000000009b90c73a26b9;
sos_loop[0].somModel.tcam_mask[7][395][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][396][0]=80'h00000000f1aad48501e0;
sos_loop[0].somModel.tcam_mask[7][396][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][397][0]=80'h00000000b50e5a5b2331;
sos_loop[0].somModel.tcam_mask[7][397][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][398][0]=80'h000000000536e70ff511;
sos_loop[0].somModel.tcam_mask[7][398][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][399][0]=80'h00000000500f137223d6;
sos_loop[0].somModel.tcam_mask[7][399][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][400][0]=80'h000000002791051b62a6;
sos_loop[0].somModel.tcam_mask[7][400][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][401][0]=80'h00000000c4eb2c045df0;
sos_loop[0].somModel.tcam_mask[7][401][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][402][0]=80'h00000000a4ad1b4e4c65;
sos_loop[0].somModel.tcam_mask[7][402][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][403][0]=80'h000000005dcd203c62ab;
sos_loop[0].somModel.tcam_mask[7][403][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][404][0]=80'h00000000bd2053fe1aa1;
sos_loop[0].somModel.tcam_mask[7][404][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][405][0]=80'h00000000dd873733eebd;
sos_loop[0].somModel.tcam_mask[7][405][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][406][0]=80'h00000000d5cc8944cc44;
sos_loop[0].somModel.tcam_mask[7][406][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][407][0]=80'h00000000df75e34c1d60;
sos_loop[0].somModel.tcam_mask[7][407][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][408][0]=80'h0000000069516c90e02b;
sos_loop[0].somModel.tcam_mask[7][408][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][409][0]=80'h00000000ba7434218648;
sos_loop[0].somModel.tcam_mask[7][409][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][410][0]=80'h0000000075995e082cc9;
sos_loop[0].somModel.tcam_mask[7][410][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][411][0]=80'h000000008f8a0618c492;
sos_loop[0].somModel.tcam_mask[7][411][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][412][0]=80'h0000000085652adefb50;
sos_loop[0].somModel.tcam_mask[7][412][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][413][0]=80'h0000000084e3bbb346a9;
sos_loop[0].somModel.tcam_mask[7][413][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][414][0]=80'h00000000ce288545ff5c;
sos_loop[0].somModel.tcam_mask[7][414][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][415][0]=80'h00000000f34840529bc7;
sos_loop[0].somModel.tcam_mask[7][415][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][416][0]=80'h0000000093b680734ca8;
sos_loop[0].somModel.tcam_mask[7][416][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][417][0]=80'h000000006d3e5930bf31;
sos_loop[0].somModel.tcam_mask[7][417][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][418][0]=80'h000000004c6bb4e13dd2;
sos_loop[0].somModel.tcam_mask[7][418][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][419][0]=80'h00000000c17e7cae146d;
sos_loop[0].somModel.tcam_mask[7][419][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][420][0]=80'h000000003a01e234f448;
sos_loop[0].somModel.tcam_mask[7][420][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][421][0]=80'h000000001f6089a70d31;
sos_loop[0].somModel.tcam_mask[7][421][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][422][0]=80'h00000000e9910acedf01;
sos_loop[0].somModel.tcam_mask[7][422][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][423][0]=80'h0000000092c1be63a45c;
sos_loop[0].somModel.tcam_mask[7][423][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][424][0]=80'h0000000077250b5545e8;
sos_loop[0].somModel.tcam_mask[7][424][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][425][0]=80'h0000000041875a4af1b4;
sos_loop[0].somModel.tcam_mask[7][425][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][426][0]=80'h000000001f7188b8f195;
sos_loop[0].somModel.tcam_mask[7][426][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][427][0]=80'h00000000e7043697f5e9;
sos_loop[0].somModel.tcam_mask[7][427][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][428][0]=80'h00000000ccb0a5325cbe;
sos_loop[0].somModel.tcam_mask[7][428][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][429][0]=80'h00000000f77c99d0ae10;
sos_loop[0].somModel.tcam_mask[7][429][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][430][0]=80'h0000000051c66267cec7;
sos_loop[0].somModel.tcam_mask[7][430][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][431][0]=80'h00000000a3eb7b517f7d;
sos_loop[0].somModel.tcam_mask[7][431][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][432][0]=80'h000000005e4b84a9a324;
sos_loop[0].somModel.tcam_mask[7][432][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][433][0]=80'h00000000263366d9a934;
sos_loop[0].somModel.tcam_mask[7][433][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][434][0]=80'h0000000035cd167e2bad;
sos_loop[0].somModel.tcam_mask[7][434][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][435][0]=80'h000000000b2c3bbf8fba;
sos_loop[0].somModel.tcam_mask[7][435][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][436][0]=80'h000000008f19a66976c7;
sos_loop[0].somModel.tcam_mask[7][436][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][437][0]=80'h00000000e0b42c35622b;
sos_loop[0].somModel.tcam_mask[7][437][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][438][0]=80'h00000000dca9a6f1782c;
sos_loop[0].somModel.tcam_mask[7][438][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][439][0]=80'h000000009a1541c274a2;
sos_loop[0].somModel.tcam_mask[7][439][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][440][0]=80'h0000000044768a38b95d;
sos_loop[0].somModel.tcam_mask[7][440][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][441][0]=80'h0000000038f48a68b142;
sos_loop[0].somModel.tcam_mask[7][441][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][442][0]=80'h000000009759c188b4fd;
sos_loop[0].somModel.tcam_mask[7][442][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][443][0]=80'h00000000a08c0f3399b6;
sos_loop[0].somModel.tcam_mask[7][443][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][444][0]=80'h00000000820dea118ef9;
sos_loop[0].somModel.tcam_mask[7][444][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][445][0]=80'h00000000786f4fec3569;
sos_loop[0].somModel.tcam_mask[7][445][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][446][0]=80'h0000000035502a9bf339;
sos_loop[0].somModel.tcam_mask[7][446][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][447][0]=80'h00000000ede032f81911;
sos_loop[0].somModel.tcam_mask[7][447][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][448][0]=80'h00000000005d2da41d57;
sos_loop[0].somModel.tcam_mask[7][448][0]=80'hffffffffff8000000000;
sos_loop[0].somModel.tcam_data[7][449][0]=80'h000000001d551e45233a;
sos_loop[0].somModel.tcam_mask[7][449][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][450][0]=80'h000000001232e7e21619;
sos_loop[0].somModel.tcam_mask[7][450][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][451][0]=80'h000000009656bf8e0b9d;
sos_loop[0].somModel.tcam_mask[7][451][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][452][0]=80'h00000000282df63c9a42;
sos_loop[0].somModel.tcam_mask[7][452][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][453][0]=80'h00000000fb8cfa3efc1a;
sos_loop[0].somModel.tcam_mask[7][453][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][454][0]=80'h00000000e202a5e04142;
sos_loop[0].somModel.tcam_mask[7][454][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][455][0]=80'h00000000ce14bd93ed55;
sos_loop[0].somModel.tcam_mask[7][455][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][456][0]=80'h000000000b29b6b75332;
sos_loop[0].somModel.tcam_mask[7][456][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][457][0]=80'h00000000a560cfe7acfc;
sos_loop[0].somModel.tcam_mask[7][457][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][458][0]=80'h0000000099c7f0448e01;
sos_loop[0].somModel.tcam_mask[7][458][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][459][0]=80'h000000001dc007e9c85a;
sos_loop[0].somModel.tcam_mask[7][459][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][460][0]=80'h00000000d5bbfcebded1;
sos_loop[0].somModel.tcam_mask[7][460][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][461][0]=80'h000000007a59ce859cc7;
sos_loop[0].somModel.tcam_mask[7][461][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][462][0]=80'h000000004ea8c5b70bda;
sos_loop[0].somModel.tcam_mask[7][462][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][463][0]=80'h0000000052f1807fc08a;
sos_loop[0].somModel.tcam_mask[7][463][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][464][0]=80'h00000000206171d9529a;
sos_loop[0].somModel.tcam_mask[7][464][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][465][0]=80'h00000000498a7ea9d6a4;
sos_loop[0].somModel.tcam_mask[7][465][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][466][0]=80'h0000000068b1d8990008;
sos_loop[0].somModel.tcam_mask[7][466][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][467][0]=80'h00000000dfdd7f5c6649;
sos_loop[0].somModel.tcam_mask[7][467][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][468][0]=80'h00000000423c83f43d47;
sos_loop[0].somModel.tcam_mask[7][468][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][469][0]=80'h0000000071daa74440c3;
sos_loop[0].somModel.tcam_mask[7][469][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][470][0]=80'h000000006b7caeb2cb69;
sos_loop[0].somModel.tcam_mask[7][470][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][471][0]=80'h000000009301716b199f;
sos_loop[0].somModel.tcam_mask[7][471][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][472][0]=80'h00000000f30c2c261355;
sos_loop[0].somModel.tcam_mask[7][472][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][473][0]=80'h00000000e1037b5789b6;
sos_loop[0].somModel.tcam_mask[7][473][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][474][0]=80'h000000004ac85c163c30;
sos_loop[0].somModel.tcam_mask[7][474][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][475][0]=80'h00000000bd2e17a3bd71;
sos_loop[0].somModel.tcam_mask[7][475][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][476][0]=80'h000000008cfbaac12a25;
sos_loop[0].somModel.tcam_mask[7][476][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][477][0]=80'h00000000e07f86b355a4;
sos_loop[0].somModel.tcam_mask[7][477][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][478][0]=80'h00000000e24b3b5f435d;
sos_loop[0].somModel.tcam_mask[7][478][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][479][0]=80'h00000000c6100a3221e3;
sos_loop[0].somModel.tcam_mask[7][479][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][480][0]=80'h00000000d601e9e5d6ac;
sos_loop[0].somModel.tcam_mask[7][480][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][481][0]=80'h00000000a2ee82f9007b;
sos_loop[0].somModel.tcam_mask[7][481][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][482][0]=80'h00000000b4baf8944204;
sos_loop[0].somModel.tcam_mask[7][482][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][483][0]=80'h0000000078c5ee1f506d;
sos_loop[0].somModel.tcam_mask[7][483][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][484][0]=80'h0000000094176a64d950;
sos_loop[0].somModel.tcam_mask[7][484][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][485][0]=80'h00000000bdc7edf2bed3;
sos_loop[0].somModel.tcam_mask[7][485][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][486][0]=80'h00000000f6141087125a;
sos_loop[0].somModel.tcam_mask[7][486][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][487][0]=80'h000000004d8a6c4bb175;
sos_loop[0].somModel.tcam_mask[7][487][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][488][0]=80'h00000000d702b7ff755e;
sos_loop[0].somModel.tcam_mask[7][488][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][489][0]=80'h0000000017ad459c4491;
sos_loop[0].somModel.tcam_mask[7][489][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][490][0]=80'h00000000becd69de0af5;
sos_loop[0].somModel.tcam_mask[7][490][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][491][0]=80'h000000006db83a09cb40;
sos_loop[0].somModel.tcam_mask[7][491][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][492][0]=80'h00000000c15a3192c54e;
sos_loop[0].somModel.tcam_mask[7][492][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][493][0]=80'h00000000372729de79a7;
sos_loop[0].somModel.tcam_mask[7][493][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][494][0]=80'h00000000b7d5a573112e;
sos_loop[0].somModel.tcam_mask[7][494][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][495][0]=80'h00000000e7598a8d64ef;
sos_loop[0].somModel.tcam_mask[7][495][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][496][0]=80'h000000004d77a8f186e8;
sos_loop[0].somModel.tcam_mask[7][496][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][497][0]=80'h00000000b3a7e8c62438;
sos_loop[0].somModel.tcam_mask[7][497][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][498][0]=80'h000000005e628e40bad8;
sos_loop[0].somModel.tcam_mask[7][498][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][499][0]=80'h000000002c6ae9566a81;
sos_loop[0].somModel.tcam_mask[7][499][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][500][0]=80'h000000007c8088a4d780;
sos_loop[0].somModel.tcam_mask[7][500][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][501][0]=80'h00000000449da718991b;
sos_loop[0].somModel.tcam_mask[7][501][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][502][0]=80'h00000000eb14915c851e;
sos_loop[0].somModel.tcam_mask[7][502][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][503][0]=80'h000000003527b3d245b5;
sos_loop[0].somModel.tcam_mask[7][503][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][504][0]=80'h0000000085d7cc131a8a;
sos_loop[0].somModel.tcam_mask[7][504][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][505][0]=80'h00000000b448dcc734b3;
sos_loop[0].somModel.tcam_mask[7][505][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][506][0]=80'h000000000463282aaf56;
sos_loop[0].somModel.tcam_mask[7][506][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][507][0]=80'h00000000e6f6fe35b667;
sos_loop[0].somModel.tcam_mask[7][507][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][508][0]=80'h0000000080c258b15826;
sos_loop[0].somModel.tcam_mask[7][508][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][509][0]=80'h00000000faac4f7283f1;
sos_loop[0].somModel.tcam_mask[7][509][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][510][0]=80'h00000000a03cce697a88;
sos_loop[0].somModel.tcam_mask[7][510][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][511][0]=80'h00000000df03c7e186d0;
sos_loop[0].somModel.tcam_mask[7][511][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][512][0]=80'h00000000c301b2ddb491;
sos_loop[0].somModel.tcam_mask[7][512][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][513][0]=80'h0000000005a553a6d946;
sos_loop[0].somModel.tcam_mask[7][513][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][514][0]=80'h00000000ec81a0ecf565;
sos_loop[0].somModel.tcam_mask[7][514][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][515][0]=80'h0000000025b7ba6c7a22;
sos_loop[0].somModel.tcam_mask[7][515][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][516][0]=80'h00000000ff62f77af68e;
sos_loop[0].somModel.tcam_mask[7][516][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][517][0]=80'h0000000090696c0e7c49;
sos_loop[0].somModel.tcam_mask[7][517][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][518][0]=80'h00000000db542752b51b;
sos_loop[0].somModel.tcam_mask[7][518][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][519][0]=80'h000000005c669d7e5719;
sos_loop[0].somModel.tcam_mask[7][519][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][520][0]=80'h0000000007869b90d6d6;
sos_loop[0].somModel.tcam_mask[7][520][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][521][0]=80'h000000006ab3f4028bc4;
sos_loop[0].somModel.tcam_mask[7][521][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][522][0]=80'h00000000faf254c81784;
sos_loop[0].somModel.tcam_mask[7][522][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][523][0]=80'h00000000e91e80ddf2b6;
sos_loop[0].somModel.tcam_mask[7][523][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][524][0]=80'h0000000012ec8002dccf;
sos_loop[0].somModel.tcam_mask[7][524][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][525][0]=80'h000000001fb66119b301;
sos_loop[0].somModel.tcam_mask[7][525][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][526][0]=80'h0000000035cfa56dca6a;
sos_loop[0].somModel.tcam_mask[7][526][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][527][0]=80'h00000000257f17287640;
sos_loop[0].somModel.tcam_mask[7][527][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][528][0]=80'h00000000e24b719e5fd5;
sos_loop[0].somModel.tcam_mask[7][528][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][529][0]=80'h000000001b6de98d63bb;
sos_loop[0].somModel.tcam_mask[7][529][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][530][0]=80'h00000000c7396a1e1d0b;
sos_loop[0].somModel.tcam_mask[7][530][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][531][0]=80'h000000007fb43ae9cd4b;
sos_loop[0].somModel.tcam_mask[7][531][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][532][0]=80'h00000000a389a8825008;
sos_loop[0].somModel.tcam_mask[7][532][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][533][0]=80'h0000000062002cc089d3;
sos_loop[0].somModel.tcam_mask[7][533][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][534][0]=80'h00000000a2fc3e097fd8;
sos_loop[0].somModel.tcam_mask[7][534][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][535][0]=80'h0000000093938f2e7bb6;
sos_loop[0].somModel.tcam_mask[7][535][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][536][0]=80'h000000004c0878c8f3c9;
sos_loop[0].somModel.tcam_mask[7][536][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][537][0]=80'h000000006dad4681d74b;
sos_loop[0].somModel.tcam_mask[7][537][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][538][0]=80'h0000000090d849afd440;
sos_loop[0].somModel.tcam_mask[7][538][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][539][0]=80'h0000000099cea5c192b2;
sos_loop[0].somModel.tcam_mask[7][539][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][540][0]=80'h00000000439a63924ef9;
sos_loop[0].somModel.tcam_mask[7][540][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][541][0]=80'h0000000022efe4c3db4e;
sos_loop[0].somModel.tcam_mask[7][541][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][542][0]=80'h00000000935f8ae1eaca;
sos_loop[0].somModel.tcam_mask[7][542][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][543][0]=80'h00000000980ce89cb3ca;
sos_loop[0].somModel.tcam_mask[7][543][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][544][0]=80'h00000000b2b1d54e6143;
sos_loop[0].somModel.tcam_mask[7][544][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][545][0]=80'h00000000985262ca09c2;
sos_loop[0].somModel.tcam_mask[7][545][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][546][0]=80'h000000001b5370c23148;
sos_loop[0].somModel.tcam_mask[7][546][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][547][0]=80'h00000000fa6e44897737;
sos_loop[0].somModel.tcam_mask[7][547][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][548][0]=80'h00000000edc347b5f551;
sos_loop[0].somModel.tcam_mask[7][548][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][549][0]=80'h00000000bbafbcb86844;
sos_loop[0].somModel.tcam_mask[7][549][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][550][0]=80'h000000007fb9ba95cb59;
sos_loop[0].somModel.tcam_mask[7][550][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][551][0]=80'h00000000be931b35ee21;
sos_loop[0].somModel.tcam_mask[7][551][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][552][0]=80'h0000000039f56d709e34;
sos_loop[0].somModel.tcam_mask[7][552][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][553][0]=80'h000000004e9dfa08200a;
sos_loop[0].somModel.tcam_mask[7][553][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][554][0]=80'h00000000820c31b21a45;
sos_loop[0].somModel.tcam_mask[7][554][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][555][0]=80'h0000000005c7809f7005;
sos_loop[0].somModel.tcam_mask[7][555][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][556][0]=80'h000000003aca0c094cca;
sos_loop[0].somModel.tcam_mask[7][556][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][557][0]=80'h00000000745ae42f60b0;
sos_loop[0].somModel.tcam_mask[7][557][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][558][0]=80'h000000009ab1034e7c6e;
sos_loop[0].somModel.tcam_mask[7][558][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][559][0]=80'h000000008b03e00b02c2;
sos_loop[0].somModel.tcam_mask[7][559][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][560][0]=80'h00000000291393c268aa;
sos_loop[0].somModel.tcam_mask[7][560][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][561][0]=80'h000000004f5dda910b46;
sos_loop[0].somModel.tcam_mask[7][561][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][562][0]=80'h000000000d702572b740;
sos_loop[0].somModel.tcam_mask[7][562][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][563][0]=80'h0000000082eb751a50eb;
sos_loop[0].somModel.tcam_mask[7][563][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][564][0]=80'h0000000069f1bf212be5;
sos_loop[0].somModel.tcam_mask[7][564][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][565][0]=80'h00000000692f8eeae2e9;
sos_loop[0].somModel.tcam_mask[7][565][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][566][0]=80'h0000000019a683169415;
sos_loop[0].somModel.tcam_mask[7][566][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][567][0]=80'h0000000093bac3e6e685;
sos_loop[0].somModel.tcam_mask[7][567][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][568][0]=80'h000000004993bee769ac;
sos_loop[0].somModel.tcam_mask[7][568][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][569][0]=80'h00000000cd7fb4cb6753;
sos_loop[0].somModel.tcam_mask[7][569][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][570][0]=80'h000000000240e7a3c36d;
sos_loop[0].somModel.tcam_mask[7][570][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[7][571][0]=80'h00000000dee7cb29be85;
sos_loop[0].somModel.tcam_mask[7][571][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][572][0]=80'h00000000992597565e42;
sos_loop[0].somModel.tcam_mask[7][572][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][573][0]=80'h000000005cf48819c736;
sos_loop[0].somModel.tcam_mask[7][573][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][574][0]=80'h0000000047abe210da7f;
sos_loop[0].somModel.tcam_mask[7][574][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][575][0]=80'h00000000f93a1757baa0;
sos_loop[0].somModel.tcam_mask[7][575][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][576][0]=80'h000000007c1ceb4afc56;
sos_loop[0].somModel.tcam_mask[7][576][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][577][0]=80'h00000000af7d256d7cc4;
sos_loop[0].somModel.tcam_mask[7][577][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][578][0]=80'h0000000056f4eacb32c7;
sos_loop[0].somModel.tcam_mask[7][578][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][579][0]=80'h00000000b0d1add53e47;
sos_loop[0].somModel.tcam_mask[7][579][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][580][0]=80'h00000000d2755cc4bd17;
sos_loop[0].somModel.tcam_mask[7][580][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][581][0]=80'h00000000a6985589f9f2;
sos_loop[0].somModel.tcam_mask[7][581][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][582][0]=80'h00000000c617a79d7ece;
sos_loop[0].somModel.tcam_mask[7][582][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][583][0]=80'h00000000ce74602fffba;
sos_loop[0].somModel.tcam_mask[7][583][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][584][0]=80'h00000000f924b4b96d61;
sos_loop[0].somModel.tcam_mask[7][584][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][585][0]=80'h000000008c0b6b9901dc;
sos_loop[0].somModel.tcam_mask[7][585][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][586][0]=80'h00000000f68af87708bf;
sos_loop[0].somModel.tcam_mask[7][586][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][587][0]=80'h0000000074fa5f30fe3f;
sos_loop[0].somModel.tcam_mask[7][587][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][588][0]=80'h000000004db8a921b1d2;
sos_loop[0].somModel.tcam_mask[7][588][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][589][0]=80'h0000000018a72f979e24;
sos_loop[0].somModel.tcam_mask[7][589][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][590][0]=80'h00000000595e18260e26;
sos_loop[0].somModel.tcam_mask[7][590][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][591][0]=80'h00000000aad2d483e822;
sos_loop[0].somModel.tcam_mask[7][591][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][592][0]=80'h00000000343913fad305;
sos_loop[0].somModel.tcam_mask[7][592][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][593][0]=80'h00000000b3d2b6c10e97;
sos_loop[0].somModel.tcam_mask[7][593][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][594][0]=80'h000000005b359f4f70b0;
sos_loop[0].somModel.tcam_mask[7][594][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][595][0]=80'h00000000910fdf65238e;
sos_loop[0].somModel.tcam_mask[7][595][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][596][0]=80'h00000000858d2a03d342;
sos_loop[0].somModel.tcam_mask[7][596][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][597][0]=80'h0000000060c0b6079327;
sos_loop[0].somModel.tcam_mask[7][597][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][598][0]=80'h00000000ac7bf03559d7;
sos_loop[0].somModel.tcam_mask[7][598][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][599][0]=80'h000000009ad2390bbe32;
sos_loop[0].somModel.tcam_mask[7][599][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][600][0]=80'h00000000fa4f7ce06718;
sos_loop[0].somModel.tcam_mask[7][600][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][601][0]=80'h00000000d16fe65ec39f;
sos_loop[0].somModel.tcam_mask[7][601][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][602][0]=80'h000000002d99e55053a9;
sos_loop[0].somModel.tcam_mask[7][602][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][603][0]=80'h000000005159029f3697;
sos_loop[0].somModel.tcam_mask[7][603][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][604][0]=80'h00000000b4b0447b5549;
sos_loop[0].somModel.tcam_mask[7][604][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][605][0]=80'h00000000377b752a37b6;
sos_loop[0].somModel.tcam_mask[7][605][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][606][0]=80'h00000000220bb11437f4;
sos_loop[0].somModel.tcam_mask[7][606][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][607][0]=80'h00000000abd69fb1204e;
sos_loop[0].somModel.tcam_mask[7][607][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][608][0]=80'h00000000eb47988d0d8b;
sos_loop[0].somModel.tcam_mask[7][608][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][609][0]=80'h00000000ca9cc767edce;
sos_loop[0].somModel.tcam_mask[7][609][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][610][0]=80'h000000003b6f42cbe0a9;
sos_loop[0].somModel.tcam_mask[7][610][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][611][0]=80'h000000001dd3fa287076;
sos_loop[0].somModel.tcam_mask[7][611][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][612][0]=80'h000000009628912dbff2;
sos_loop[0].somModel.tcam_mask[7][612][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][613][0]=80'h0000000089a7951bea35;
sos_loop[0].somModel.tcam_mask[7][613][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][614][0]=80'h00000000c7b2ff90ab75;
sos_loop[0].somModel.tcam_mask[7][614][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][615][0]=80'h000000007ec37d3f35d1;
sos_loop[0].somModel.tcam_mask[7][615][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][616][0]=80'h00000000486d45350ba4;
sos_loop[0].somModel.tcam_mask[7][616][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][617][0]=80'h00000000f7c78a4aeffd;
sos_loop[0].somModel.tcam_mask[7][617][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][618][0]=80'h00000000ea7f3c4470a0;
sos_loop[0].somModel.tcam_mask[7][618][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][619][0]=80'h0000000095398bca46db;
sos_loop[0].somModel.tcam_mask[7][619][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][620][0]=80'h0000000002a21d269ef9;
sos_loop[0].somModel.tcam_mask[7][620][0]=80'hfffffffffc0000000000;
sos_loop[0].somModel.tcam_data[7][621][0]=80'h000000005ff142432afa;
sos_loop[0].somModel.tcam_mask[7][621][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][622][0]=80'h000000008d346fc65e2b;
sos_loop[0].somModel.tcam_mask[7][622][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][623][0]=80'h000000001a6584f50556;
sos_loop[0].somModel.tcam_mask[7][623][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][624][0]=80'h0000000008386da1029f;
sos_loop[0].somModel.tcam_mask[7][624][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][625][0]=80'h00000000db56c981ece6;
sos_loop[0].somModel.tcam_mask[7][625][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][626][0]=80'h00000000cfe8af38f522;
sos_loop[0].somModel.tcam_mask[7][626][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][627][0]=80'h000000008e919d8a745b;
sos_loop[0].somModel.tcam_mask[7][627][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][628][0]=80'h00000000543818958c78;
sos_loop[0].somModel.tcam_mask[7][628][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][629][0]=80'h00000000a8b931f97188;
sos_loop[0].somModel.tcam_mask[7][629][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][630][0]=80'h000000007dee0d849922;
sos_loop[0].somModel.tcam_mask[7][630][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][631][0]=80'h000000001017ca8a2953;
sos_loop[0].somModel.tcam_mask[7][631][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][632][0]=80'h000000007ed9cae24403;
sos_loop[0].somModel.tcam_mask[7][632][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][633][0]=80'h00000000ea187ed4d55a;
sos_loop[0].somModel.tcam_mask[7][633][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][634][0]=80'h000000002e76e28270f1;
sos_loop[0].somModel.tcam_mask[7][634][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][635][0]=80'h00000000f1980343333f;
sos_loop[0].somModel.tcam_mask[7][635][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][636][0]=80'h000000008de1c963c062;
sos_loop[0].somModel.tcam_mask[7][636][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][637][0]=80'h000000003fd86ea44501;
sos_loop[0].somModel.tcam_mask[7][637][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][638][0]=80'h00000000dc791a00bf2c;
sos_loop[0].somModel.tcam_mask[7][638][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][639][0]=80'h0000000076fd772b3105;
sos_loop[0].somModel.tcam_mask[7][639][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][640][0]=80'h000000009137a6d429b2;
sos_loop[0].somModel.tcam_mask[7][640][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][641][0]=80'h0000000049d4cbef7ccc;
sos_loop[0].somModel.tcam_mask[7][641][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][642][0]=80'h000000008051f12b529f;
sos_loop[0].somModel.tcam_mask[7][642][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][643][0]=80'h0000000008d6aa657a5e;
sos_loop[0].somModel.tcam_mask[7][643][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][644][0]=80'h0000000044bafb829ee6;
sos_loop[0].somModel.tcam_mask[7][644][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][645][0]=80'h00000000e55061ccc7b7;
sos_loop[0].somModel.tcam_mask[7][645][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][646][0]=80'h00000000d75970bd3bb0;
sos_loop[0].somModel.tcam_mask[7][646][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][647][0]=80'h000000004811729ba385;
sos_loop[0].somModel.tcam_mask[7][647][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][648][0]=80'h00000000c0501fd955df;
sos_loop[0].somModel.tcam_mask[7][648][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][649][0]=80'h00000000659c29b06d69;
sos_loop[0].somModel.tcam_mask[7][649][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][650][0]=80'h000000006aec373261a3;
sos_loop[0].somModel.tcam_mask[7][650][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][651][0]=80'h00000000c25cd90f5dab;
sos_loop[0].somModel.tcam_mask[7][651][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][652][0]=80'h00000000cee3230bfef6;
sos_loop[0].somModel.tcam_mask[7][652][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][653][0]=80'h000000007bde198a992f;
sos_loop[0].somModel.tcam_mask[7][653][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][654][0]=80'h000000007cd4d9587ccb;
sos_loop[0].somModel.tcam_mask[7][654][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][655][0]=80'h000000005cee7e94dd42;
sos_loop[0].somModel.tcam_mask[7][655][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][656][0]=80'h000000000c7f2c96b613;
sos_loop[0].somModel.tcam_mask[7][656][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][657][0]=80'h00000000f2de9d0bdde4;
sos_loop[0].somModel.tcam_mask[7][657][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][658][0]=80'h00000000b80342294761;
sos_loop[0].somModel.tcam_mask[7][658][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][659][0]=80'h00000000ef05f9051dde;
sos_loop[0].somModel.tcam_mask[7][659][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][660][0]=80'h00000000089d9864b0f7;
sos_loop[0].somModel.tcam_mask[7][660][0]=80'hfffffffff00000000000;
sos_loop[0].somModel.tcam_data[7][661][0]=80'h00000000f84ebc6b5933;
sos_loop[0].somModel.tcam_mask[7][661][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][662][0]=80'h0000000099c7ebd6ef11;
sos_loop[0].somModel.tcam_mask[7][662][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][663][0]=80'h00000000a5cfc726453c;
sos_loop[0].somModel.tcam_mask[7][663][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][664][0]=80'h000000008e33ccc43905;
sos_loop[0].somModel.tcam_mask[7][664][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][665][0]=80'h0000000061dbc393f8b8;
sos_loop[0].somModel.tcam_mask[7][665][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][666][0]=80'h00000000b5776eb8e40c;
sos_loop[0].somModel.tcam_mask[7][666][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][667][0]=80'h00000000c56f02fbb8af;
sos_loop[0].somModel.tcam_mask[7][667][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][668][0]=80'h00000000f06ac89a6e2e;
sos_loop[0].somModel.tcam_mask[7][668][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][669][0]=80'h000000004d46ea5704c7;
sos_loop[0].somModel.tcam_mask[7][669][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][670][0]=80'h00000000018a0d2ab536;
sos_loop[0].somModel.tcam_mask[7][670][0]=80'hfffffffffe0000000000;
sos_loop[0].somModel.tcam_data[7][671][0]=80'h00000000de24ea9c8559;
sos_loop[0].somModel.tcam_mask[7][671][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][672][0]=80'h00000000117c2dcb8a3f;
sos_loop[0].somModel.tcam_mask[7][672][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][673][0]=80'h00000000042c5800a198;
sos_loop[0].somModel.tcam_mask[7][673][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][674][0]=80'h00000000c866641162c8;
sos_loop[0].somModel.tcam_mask[7][674][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][675][0]=80'h00000000c59ce2a178ef;
sos_loop[0].somModel.tcam_mask[7][675][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][676][0]=80'h0000000091b9a88b2186;
sos_loop[0].somModel.tcam_mask[7][676][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][677][0]=80'h00000000baaaa92f9330;
sos_loop[0].somModel.tcam_mask[7][677][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][678][0]=80'h00000000899bc4d45fed;
sos_loop[0].somModel.tcam_mask[7][678][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][679][0]=80'h0000000031aba86c07cd;
sos_loop[0].somModel.tcam_mask[7][679][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][680][0]=80'h00000000c4984e56b9a3;
sos_loop[0].somModel.tcam_mask[7][680][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][681][0]=80'h000000001b2cb5378bd2;
sos_loop[0].somModel.tcam_mask[7][681][0]=80'hffffffffe00000000000;
sos_loop[0].somModel.tcam_data[7][682][0]=80'h00000000ff120ca68f9a;
sos_loop[0].somModel.tcam_mask[7][682][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][683][0]=80'h00000000a835dfd4a64e;
sos_loop[0].somModel.tcam_mask[7][683][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][684][0]=80'h00000000cc35683c57dc;
sos_loop[0].somModel.tcam_mask[7][684][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][685][0]=80'h00000000a5c1099a0ccc;
sos_loop[0].somModel.tcam_mask[7][685][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][686][0]=80'h00000000efd95c4e5fe9;
sos_loop[0].somModel.tcam_mask[7][686][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][687][0]=80'h000000007c76d25796aa;
sos_loop[0].somModel.tcam_mask[7][687][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][688][0]=80'h0000000007b60730923d;
sos_loop[0].somModel.tcam_mask[7][688][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][689][0]=80'h0000000007373b8b8f3c;
sos_loop[0].somModel.tcam_mask[7][689][0]=80'hfffffffff80000000000;
sos_loop[0].somModel.tcam_data[7][690][0]=80'h0000000037e56c799b77;
sos_loop[0].somModel.tcam_mask[7][690][0]=80'hffffffffc00000000000;
sos_loop[0].somModel.tcam_data[7][691][0]=80'h0000000064aeec7ab84c;
sos_loop[0].somModel.tcam_mask[7][691][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][692][0]=80'h00000000dc1814387312;
sos_loop[0].somModel.tcam_mask[7][692][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][693][0]=80'h00000000dd2835b8c4f9;
sos_loop[0].somModel.tcam_mask[7][693][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][694][0]=80'h000000005af2eb552cca;
sos_loop[0].somModel.tcam_mask[7][694][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][695][0]=80'h00000000446b9299fa74;
sos_loop[0].somModel.tcam_mask[7][695][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][696][0]=80'h0000000086928cf64fc6;
sos_loop[0].somModel.tcam_mask[7][696][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][697][0]=80'h00000000c4fdc019c61f;
sos_loop[0].somModel.tcam_mask[7][697][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][698][0]=80'h00000000882f97bb161f;
sos_loop[0].somModel.tcam_mask[7][698][0]=80'hffffffff000000000000;
sos_loop[0].somModel.tcam_data[7][699][0]=80'h000000004ed606f4518d;
sos_loop[0].somModel.tcam_mask[7][699][0]=80'hffffffff800000000000;
sos_loop[0].somModel.tcam_data[7][700][0]=80'h00000000bd46a3aa3c15;
sos_loop[0].somModel.tcam_mask[7][700][0]=80'hffffffff000000000000;
sos_loop[0].somModel.sram_dat[7][0][0]=96'hdeadbf;
sos_loop[0].somModel.sram_ptr[7][0]=939;
sos_loop[0].somModel.sram_dat[7][1][0]=96'h6814;
sos_loop[0].somModel.sram_ptr[7][1]=3;
sos_loop[0].somModel.sram_dat[7][2][0]=96'hc070;
sos_loop[0].somModel.sram_ptr[7][2]=3;
sos_loop[0].somModel.sram_dat[7][3][0]=96'h9740;
sos_loop[0].somModel.sram_ptr[7][3]=3;
sos_loop[0].somModel.sram_dat[7][4][0]=96'hc6fc;
sos_loop[0].somModel.sram_ptr[7][4]=3;
sos_loop[0].somModel.sram_dat[7][5][0]=96'h123a;
sos_loop[0].somModel.sram_ptr[7][5]=3;
sos_loop[0].somModel.sram_dat[7][6][0]=96'h7780;
sos_loop[0].somModel.sram_ptr[7][6]=3;
sos_loop[0].somModel.sram_dat[7][7][0]=96'ha3a1;
sos_loop[0].somModel.sram_ptr[7][7]=3;
sos_loop[0].somModel.sram_dat[7][8][0]=96'h3259;
sos_loop[0].somModel.sram_ptr[7][8]=3;
sos_loop[0].somModel.sram_dat[7][9][0]=96'hb3e9;
sos_loop[0].somModel.sram_ptr[7][9]=3;
sos_loop[0].somModel.sram_dat[7][10][0]=96'h6bec;
sos_loop[0].somModel.sram_ptr[7][10]=3;
sos_loop[0].somModel.sram_dat[7][11][0]=96'h3843;
sos_loop[0].somModel.sram_ptr[7][11]=3;
sos_loop[0].somModel.sram_dat[7][12][0]=96'h89af;
sos_loop[0].somModel.sram_ptr[7][12]=3;
sos_loop[0].somModel.sram_dat[7][13][0]=96'h8c78;
sos_loop[0].somModel.sram_ptr[7][13]=3;
sos_loop[0].somModel.sram_dat[7][14][0]=96'h18e7;
sos_loop[0].somModel.sram_ptr[7][14]=3;
sos_loop[0].somModel.sram_dat[7][15][0]=96'h75ae;
sos_loop[0].somModel.sram_ptr[7][15]=3;
sos_loop[0].somModel.sram_dat[7][16][0]=96'h80c5;
sos_loop[0].somModel.sram_ptr[7][16]=3;
sos_loop[0].somModel.sram_dat[7][17][0]=96'h9a32;
sos_loop[0].somModel.sram_ptr[7][17]=3;
sos_loop[0].somModel.sram_dat[7][18][0]=96'he7a9;
sos_loop[0].somModel.sram_ptr[7][18]=3;
sos_loop[0].somModel.sram_dat[7][19][0]=96'hebf7;
sos_loop[0].somModel.sram_ptr[7][19]=3;
sos_loop[0].somModel.sram_dat[7][20][0]=96'hcd9a;
sos_loop[0].somModel.sram_ptr[7][20]=3;
sos_loop[0].somModel.sram_dat[7][21][0]=96'h2365;
sos_loop[0].somModel.sram_ptr[7][21]=3;
sos_loop[0].somModel.sram_dat[7][22][0]=96'h9688;
sos_loop[0].somModel.sram_ptr[7][22]=3;
sos_loop[0].somModel.sram_dat[7][23][0]=96'he859;
sos_loop[0].somModel.sram_ptr[7][23]=3;
sos_loop[0].somModel.sram_dat[7][24][0]=96'hb77b;
sos_loop[0].somModel.sram_ptr[7][24]=3;
sos_loop[0].somModel.sram_dat[7][25][0]=96'h2430;
sos_loop[0].somModel.sram_ptr[7][25]=3;
sos_loop[0].somModel.sram_dat[7][26][0]=96'hcb20;
sos_loop[0].somModel.sram_ptr[7][26]=3;
sos_loop[0].somModel.sram_dat[7][27][0]=96'ha1e3;
sos_loop[0].somModel.sram_ptr[7][27]=3;
sos_loop[0].somModel.sram_dat[7][28][0]=96'hacc;
sos_loop[0].somModel.sram_ptr[7][28]=3;
sos_loop[0].somModel.sram_dat[7][29][0]=96'heb72;
sos_loop[0].somModel.sram_ptr[7][29]=3;
sos_loop[0].somModel.sram_dat[7][30][0]=96'hf78;
sos_loop[0].somModel.sram_ptr[7][30]=3;
sos_loop[0].somModel.sram_dat[7][31][0]=96'h7d85;
sos_loop[0].somModel.sram_ptr[7][31]=3;
sos_loop[0].somModel.sram_dat[7][32][0]=96'hd586;
sos_loop[0].somModel.sram_ptr[7][32]=3;
sos_loop[0].somModel.sram_dat[7][33][0]=96'h7dab;
sos_loop[0].somModel.sram_ptr[7][33]=3;
sos_loop[0].somModel.sram_dat[7][34][0]=96'hcb04;
sos_loop[0].somModel.sram_ptr[7][34]=3;
sos_loop[0].somModel.sram_dat[7][35][0]=96'h9cbc;
sos_loop[0].somModel.sram_ptr[7][35]=3;
sos_loop[0].somModel.sram_dat[7][36][0]=96'he211;
sos_loop[0].somModel.sram_ptr[7][36]=3;
sos_loop[0].somModel.sram_dat[7][37][0]=96'hb146;
sos_loop[0].somModel.sram_ptr[7][37]=3;
sos_loop[0].somModel.sram_dat[7][38][0]=96'h4e87;
sos_loop[0].somModel.sram_ptr[7][38]=3;
sos_loop[0].somModel.sram_dat[7][39][0]=96'h597c;
sos_loop[0].somModel.sram_ptr[7][39]=3;
sos_loop[0].somModel.sram_dat[7][40][0]=96'h3e12;
sos_loop[0].somModel.sram_ptr[7][40]=3;
sos_loop[0].somModel.sram_dat[7][41][0]=96'h9949;
sos_loop[0].somModel.sram_ptr[7][41]=3;
sos_loop[0].somModel.sram_dat[7][42][0]=96'h94fa;
sos_loop[0].somModel.sram_ptr[7][42]=3;
sos_loop[0].somModel.sram_dat[7][43][0]=96'hcdb2;
sos_loop[0].somModel.sram_ptr[7][43]=3;
sos_loop[0].somModel.sram_dat[7][44][0]=96'hfe66;
sos_loop[0].somModel.sram_ptr[7][44]=3;
sos_loop[0].somModel.sram_dat[7][45][0]=96'hc0c2;
sos_loop[0].somModel.sram_ptr[7][45]=3;
sos_loop[0].somModel.sram_dat[7][46][0]=96'hf232;
sos_loop[0].somModel.sram_ptr[7][46]=3;
sos_loop[0].somModel.sram_dat[7][47][0]=96'ha7be;
sos_loop[0].somModel.sram_ptr[7][47]=3;
sos_loop[0].somModel.sram_dat[7][48][0]=96'hfcd;
sos_loop[0].somModel.sram_ptr[7][48]=3;
sos_loop[0].somModel.sram_dat[7][49][0]=96'hb422;
sos_loop[0].somModel.sram_ptr[7][49]=3;
sos_loop[0].somModel.sram_dat[7][50][0]=96'hd35e;
sos_loop[0].somModel.sram_ptr[7][50]=3;
sos_loop[0].somModel.sram_dat[7][51][0]=96'ha927;
sos_loop[0].somModel.sram_ptr[7][51]=3;
sos_loop[0].somModel.sram_dat[7][52][0]=96'hb0b8;
sos_loop[0].somModel.sram_ptr[7][52]=3;
sos_loop[0].somModel.sram_dat[7][53][0]=96'h6f6b;
sos_loop[0].somModel.sram_ptr[7][53]=3;
sos_loop[0].somModel.sram_dat[7][54][0]=96'hbd1d;
sos_loop[0].somModel.sram_ptr[7][54]=3;
sos_loop[0].somModel.sram_dat[7][55][0]=96'h981d;
sos_loop[0].somModel.sram_ptr[7][55]=3;
sos_loop[0].somModel.sram_dat[7][56][0]=96'hafd;
sos_loop[0].somModel.sram_ptr[7][56]=3;
sos_loop[0].somModel.sram_dat[7][57][0]=96'hdd25;
sos_loop[0].somModel.sram_ptr[7][57]=3;
sos_loop[0].somModel.sram_dat[7][58][0]=96'h6dac;
sos_loop[0].somModel.sram_ptr[7][58]=3;
sos_loop[0].somModel.sram_dat[7][59][0]=96'h25d5;
sos_loop[0].somModel.sram_ptr[7][59]=3;
sos_loop[0].somModel.sram_dat[7][60][0]=96'h5737;
sos_loop[0].somModel.sram_ptr[7][60]=3;
sos_loop[0].somModel.sram_dat[7][61][0]=96'h964f;
sos_loop[0].somModel.sram_ptr[7][61]=3;
sos_loop[0].somModel.sram_dat[7][62][0]=96'hee96;
sos_loop[0].somModel.sram_ptr[7][62]=3;
sos_loop[0].somModel.sram_dat[7][63][0]=96'h8464;
sos_loop[0].somModel.sram_ptr[7][63]=3;
sos_loop[0].somModel.sram_dat[7][64][0]=96'hbe76;
sos_loop[0].somModel.sram_ptr[7][64]=3;
sos_loop[0].somModel.sram_dat[7][65][0]=96'h5a21;
sos_loop[0].somModel.sram_ptr[7][65]=3;
sos_loop[0].somModel.sram_dat[7][66][0]=96'h550d;
sos_loop[0].somModel.sram_ptr[7][66]=3;
sos_loop[0].somModel.sram_dat[7][67][0]=96'hebb4;
sos_loop[0].somModel.sram_ptr[7][67]=3;
sos_loop[0].somModel.sram_dat[7][68][0]=96'hcc55;
sos_loop[0].somModel.sram_ptr[7][68]=3;
sos_loop[0].somModel.sram_dat[7][69][0]=96'h7a15;
sos_loop[0].somModel.sram_ptr[7][69]=3;
sos_loop[0].somModel.sram_dat[7][70][0]=96'hd887;
sos_loop[0].somModel.sram_ptr[7][70]=3;
sos_loop[0].somModel.sram_dat[7][71][0]=96'h6379;
sos_loop[0].somModel.sram_ptr[7][71]=3;
sos_loop[0].somModel.sram_dat[7][72][0]=96'h843c;
sos_loop[0].somModel.sram_ptr[7][72]=3;
sos_loop[0].somModel.sram_dat[7][73][0]=96'h353c;
sos_loop[0].somModel.sram_ptr[7][73]=3;
sos_loop[0].somModel.sram_dat[7][74][0]=96'h43e1;
sos_loop[0].somModel.sram_ptr[7][74]=3;
sos_loop[0].somModel.sram_dat[7][75][0]=96'h9c19;
sos_loop[0].somModel.sram_ptr[7][75]=3;
sos_loop[0].somModel.sram_dat[7][76][0]=96'hcd0b;
sos_loop[0].somModel.sram_ptr[7][76]=3;
sos_loop[0].somModel.sram_dat[7][77][0]=96'h5254;
sos_loop[0].somModel.sram_ptr[7][77]=3;
sos_loop[0].somModel.sram_dat[7][78][0]=96'hd8e8;
sos_loop[0].somModel.sram_ptr[7][78]=3;
sos_loop[0].somModel.sram_dat[7][79][0]=96'he7a6;
sos_loop[0].somModel.sram_ptr[7][79]=3;
sos_loop[0].somModel.sram_dat[7][80][0]=96'ha32f;
sos_loop[0].somModel.sram_ptr[7][80]=3;
sos_loop[0].somModel.sram_dat[7][81][0]=96'hfb8d;
sos_loop[0].somModel.sram_ptr[7][81]=3;
sos_loop[0].somModel.sram_dat[7][82][0]=96'h39f9;
sos_loop[0].somModel.sram_ptr[7][82]=3;
sos_loop[0].somModel.sram_dat[7][83][0]=96'h7d79;
sos_loop[0].somModel.sram_ptr[7][83]=3;
sos_loop[0].somModel.sram_dat[7][84][0]=96'hb263;
sos_loop[0].somModel.sram_ptr[7][84]=3;
sos_loop[0].somModel.sram_dat[7][85][0]=96'hb28d;
sos_loop[0].somModel.sram_ptr[7][85]=3;
sos_loop[0].somModel.sram_dat[7][86][0]=96'h5639;
sos_loop[0].somModel.sram_ptr[7][86]=3;
sos_loop[0].somModel.sram_dat[7][87][0]=96'h2011;
sos_loop[0].somModel.sram_ptr[7][87]=3;
sos_loop[0].somModel.sram_dat[7][88][0]=96'hbf31;
sos_loop[0].somModel.sram_ptr[7][88]=3;
sos_loop[0].somModel.sram_dat[7][89][0]=96'h902b;
sos_loop[0].somModel.sram_ptr[7][89]=3;
sos_loop[0].somModel.sram_dat[7][90][0]=96'h889d;
sos_loop[0].somModel.sram_ptr[7][90]=3;
sos_loop[0].somModel.sram_dat[7][91][0]=96'h1e7e;
sos_loop[0].somModel.sram_ptr[7][91]=3;
sos_loop[0].somModel.sram_dat[7][92][0]=96'h66b7;
sos_loop[0].somModel.sram_ptr[7][92]=3;
sos_loop[0].somModel.sram_dat[7][93][0]=96'he7a4;
sos_loop[0].somModel.sram_ptr[7][93]=3;
sos_loop[0].somModel.sram_dat[7][94][0]=96'hf191;
sos_loop[0].somModel.sram_ptr[7][94]=3;
sos_loop[0].somModel.sram_dat[7][95][0]=96'ha000;
sos_loop[0].somModel.sram_ptr[7][95]=3;
sos_loop[0].somModel.sram_dat[7][96][0]=96'h304f;
sos_loop[0].somModel.sram_ptr[7][96]=3;
sos_loop[0].somModel.sram_dat[7][97][0]=96'hcc62;
sos_loop[0].somModel.sram_ptr[7][97]=3;
sos_loop[0].somModel.sram_dat[7][98][0]=96'h42cd;
sos_loop[0].somModel.sram_ptr[7][98]=3;
sos_loop[0].somModel.sram_dat[7][99][0]=96'hb26a;
sos_loop[0].somModel.sram_ptr[7][99]=3;
sos_loop[0].somModel.sram_dat[7][100][0]=96'hc7be;
sos_loop[0].somModel.sram_ptr[7][100]=3;
sos_loop[0].somModel.sram_dat[7][101][0]=96'hb1b8;
sos_loop[0].somModel.sram_ptr[7][101]=3;
sos_loop[0].somModel.sram_dat[7][102][0]=96'hfac7;
sos_loop[0].somModel.sram_ptr[7][102]=3;
sos_loop[0].somModel.sram_dat[7][103][0]=96'h22e7;
sos_loop[0].somModel.sram_ptr[7][103]=3;
sos_loop[0].somModel.sram_dat[7][104][0]=96'h85e;
sos_loop[0].somModel.sram_ptr[7][104]=3;
sos_loop[0].somModel.sram_dat[7][105][0]=96'h6156;
sos_loop[0].somModel.sram_ptr[7][105]=3;
sos_loop[0].somModel.sram_dat[7][106][0]=96'h4e18;
sos_loop[0].somModel.sram_ptr[7][106]=3;
sos_loop[0].somModel.sram_dat[7][107][0]=96'h8df4;
sos_loop[0].somModel.sram_ptr[7][107]=3;
sos_loop[0].somModel.sram_dat[7][108][0]=96'hc184;
sos_loop[0].somModel.sram_ptr[7][108]=3;
sos_loop[0].somModel.sram_dat[7][109][0]=96'h24f9;
sos_loop[0].somModel.sram_ptr[7][109]=3;
sos_loop[0].somModel.sram_dat[7][110][0]=96'h55a9;
sos_loop[0].somModel.sram_ptr[7][110]=3;
sos_loop[0].somModel.sram_dat[7][111][0]=96'h7d2c;
sos_loop[0].somModel.sram_ptr[7][111]=3;
sos_loop[0].somModel.sram_dat[7][112][0]=96'h8b7b;
sos_loop[0].somModel.sram_ptr[7][112]=3;
sos_loop[0].somModel.sram_dat[7][113][0]=96'h6e62;
sos_loop[0].somModel.sram_ptr[7][113]=3;
sos_loop[0].somModel.sram_dat[7][114][0]=96'haa01;
sos_loop[0].somModel.sram_ptr[7][114]=3;
sos_loop[0].somModel.sram_dat[7][115][0]=96'hb523;
sos_loop[0].somModel.sram_ptr[7][115]=3;
sos_loop[0].somModel.sram_dat[7][116][0]=96'h9dba;
sos_loop[0].somModel.sram_ptr[7][116]=3;
sos_loop[0].somModel.sram_dat[7][117][0]=96'hc4e7;
sos_loop[0].somModel.sram_ptr[7][117]=3;
sos_loop[0].somModel.sram_dat[7][118][0]=96'hdf70;
sos_loop[0].somModel.sram_ptr[7][118]=3;
sos_loop[0].somModel.sram_dat[7][119][0]=96'ha6b;
sos_loop[0].somModel.sram_ptr[7][119]=3;
sos_loop[0].somModel.sram_dat[7][120][0]=96'h3efb;
sos_loop[0].somModel.sram_ptr[7][120]=3;
sos_loop[0].somModel.sram_dat[7][121][0]=96'hc13b;
sos_loop[0].somModel.sram_ptr[7][121]=3;
sos_loop[0].somModel.sram_dat[7][122][0]=96'hdd53;
sos_loop[0].somModel.sram_ptr[7][122]=3;
sos_loop[0].somModel.sram_dat[7][123][0]=96'hdc42;
sos_loop[0].somModel.sram_ptr[7][123]=3;
sos_loop[0].somModel.sram_dat[7][124][0]=96'hd019;
sos_loop[0].somModel.sram_ptr[7][124]=3;
sos_loop[0].somModel.sram_dat[7][125][0]=96'h4ac7;
sos_loop[0].somModel.sram_ptr[7][125]=3;
sos_loop[0].somModel.sram_dat[7][126][0]=96'h1c65;
sos_loop[0].somModel.sram_ptr[7][126]=3;
sos_loop[0].somModel.sram_dat[7][127][0]=96'hc12e;
sos_loop[0].somModel.sram_ptr[7][127]=3;
sos_loop[0].somModel.sram_dat[7][128][0]=96'h6cc2;
sos_loop[0].somModel.sram_ptr[7][128]=3;
sos_loop[0].somModel.sram_dat[7][129][0]=96'h1979;
sos_loop[0].somModel.sram_ptr[7][129]=3;
sos_loop[0].somModel.sram_dat[7][130][0]=96'h3003;
sos_loop[0].somModel.sram_ptr[7][130]=3;
sos_loop[0].somModel.sram_dat[7][131][0]=96'he7fc;
sos_loop[0].somModel.sram_ptr[7][131]=3;
sos_loop[0].somModel.sram_dat[7][132][0]=96'hb67b;
sos_loop[0].somModel.sram_ptr[7][132]=3;
sos_loop[0].somModel.sram_dat[7][133][0]=96'hd14d;
sos_loop[0].somModel.sram_ptr[7][133]=3;
sos_loop[0].somModel.sram_dat[7][134][0]=96'h8684;
sos_loop[0].somModel.sram_ptr[7][134]=3;
sos_loop[0].somModel.sram_dat[7][135][0]=96'h6940;
sos_loop[0].somModel.sram_ptr[7][135]=3;
sos_loop[0].somModel.sram_dat[7][136][0]=96'h34fd;
sos_loop[0].somModel.sram_ptr[7][136]=3;
sos_loop[0].somModel.sram_dat[7][137][0]=96'h89e2;
sos_loop[0].somModel.sram_ptr[7][137]=3;
sos_loop[0].somModel.sram_dat[7][138][0]=96'hda12;
sos_loop[0].somModel.sram_ptr[7][138]=3;
sos_loop[0].somModel.sram_dat[7][139][0]=96'h864;
sos_loop[0].somModel.sram_ptr[7][139]=3;
sos_loop[0].somModel.sram_dat[7][140][0]=96'hb1ee;
sos_loop[0].somModel.sram_ptr[7][140]=3;
sos_loop[0].somModel.sram_dat[7][141][0]=96'hb1e4;
sos_loop[0].somModel.sram_ptr[7][141]=3;
sos_loop[0].somModel.sram_dat[7][142][0]=96'hcc72;
sos_loop[0].somModel.sram_ptr[7][142]=3;
sos_loop[0].somModel.sram_dat[7][143][0]=96'hbe14;
sos_loop[0].somModel.sram_ptr[7][143]=3;
sos_loop[0].somModel.sram_dat[7][144][0]=96'hcda4;
sos_loop[0].somModel.sram_ptr[7][144]=3;
sos_loop[0].somModel.sram_dat[7][145][0]=96'h40c1;
sos_loop[0].somModel.sram_ptr[7][145]=3;
sos_loop[0].somModel.sram_dat[7][146][0]=96'h5d6d;
sos_loop[0].somModel.sram_ptr[7][146]=3;
sos_loop[0].somModel.sram_dat[7][147][0]=96'h4fc3;
sos_loop[0].somModel.sram_ptr[7][147]=3;
sos_loop[0].somModel.sram_dat[7][148][0]=96'hc62b;
sos_loop[0].somModel.sram_ptr[7][148]=3;
sos_loop[0].somModel.sram_dat[7][149][0]=96'hf641;
sos_loop[0].somModel.sram_ptr[7][149]=3;
sos_loop[0].somModel.sram_dat[7][150][0]=96'hcef3;
sos_loop[0].somModel.sram_ptr[7][150]=3;
sos_loop[0].somModel.sram_dat[7][151][0]=96'h585;
sos_loop[0].somModel.sram_ptr[7][151]=3;
sos_loop[0].somModel.sram_dat[7][152][0]=96'h58e;
sos_loop[0].somModel.sram_ptr[7][152]=3;
sos_loop[0].somModel.sram_dat[7][153][0]=96'h8895;
sos_loop[0].somModel.sram_ptr[7][153]=3;
sos_loop[0].somModel.sram_dat[7][154][0]=96'h8e73;
sos_loop[0].somModel.sram_ptr[7][154]=3;
sos_loop[0].somModel.sram_dat[7][155][0]=96'hbc7d;
sos_loop[0].somModel.sram_ptr[7][155]=3;
sos_loop[0].somModel.sram_dat[7][156][0]=96'hd48;
sos_loop[0].somModel.sram_ptr[7][156]=3;
sos_loop[0].somModel.sram_dat[7][157][0]=96'hde40;
sos_loop[0].somModel.sram_ptr[7][157]=3;
sos_loop[0].somModel.sram_dat[7][158][0]=96'hc40;
sos_loop[0].somModel.sram_ptr[7][158]=3;
sos_loop[0].somModel.sram_dat[7][159][0]=96'h200d;
sos_loop[0].somModel.sram_ptr[7][159]=3;
sos_loop[0].somModel.sram_dat[7][160][0]=96'h1ac3;
sos_loop[0].somModel.sram_ptr[7][160]=3;
sos_loop[0].somModel.sram_dat[7][161][0]=96'h7006;
sos_loop[0].somModel.sram_ptr[7][161]=3;
sos_loop[0].somModel.sram_dat[7][162][0]=96'hbc2d;
sos_loop[0].somModel.sram_ptr[7][162]=3;
sos_loop[0].somModel.sram_dat[7][163][0]=96'hda27;
sos_loop[0].somModel.sram_ptr[7][163]=3;
sos_loop[0].somModel.sram_dat[7][164][0]=96'he8d9;
sos_loop[0].somModel.sram_ptr[7][164]=3;
sos_loop[0].somModel.sram_dat[7][165][0]=96'hcf50;
sos_loop[0].somModel.sram_ptr[7][165]=3;
sos_loop[0].somModel.sram_dat[7][166][0]=96'h53d6;
sos_loop[0].somModel.sram_ptr[7][166]=3;
sos_loop[0].somModel.sram_dat[7][167][0]=96'h8515;
sos_loop[0].somModel.sram_ptr[7][167]=3;
sos_loop[0].somModel.sram_dat[7][168][0]=96'h3f78;
sos_loop[0].somModel.sram_ptr[7][168]=3;
sos_loop[0].somModel.sram_dat[7][169][0]=96'hf457;
sos_loop[0].somModel.sram_ptr[7][169]=3;
sos_loop[0].somModel.sram_dat[7][170][0]=96'h44bc;
sos_loop[0].somModel.sram_ptr[7][170]=3;
sos_loop[0].somModel.sram_dat[7][171][0]=96'hea98;
sos_loop[0].somModel.sram_ptr[7][171]=3;
sos_loop[0].somModel.sram_dat[7][172][0]=96'h8e43;
sos_loop[0].somModel.sram_ptr[7][172]=3;
sos_loop[0].somModel.sram_dat[7][173][0]=96'h2164;
sos_loop[0].somModel.sram_ptr[7][173]=3;
sos_loop[0].somModel.sram_dat[7][174][0]=96'h3319;
sos_loop[0].somModel.sram_ptr[7][174]=3;
sos_loop[0].somModel.sram_dat[7][175][0]=96'ha7d4;
sos_loop[0].somModel.sram_ptr[7][175]=3;
sos_loop[0].somModel.sram_dat[7][176][0]=96'h32a8;
sos_loop[0].somModel.sram_ptr[7][176]=3;
sos_loop[0].somModel.sram_dat[7][177][0]=96'he83b;
sos_loop[0].somModel.sram_ptr[7][177]=3;
sos_loop[0].somModel.sram_dat[7][178][0]=96'h1fb9;
sos_loop[0].somModel.sram_ptr[7][178]=3;
sos_loop[0].somModel.sram_dat[7][179][0]=96'h97e4;
sos_loop[0].somModel.sram_ptr[7][179]=3;
sos_loop[0].somModel.sram_dat[7][180][0]=96'hc832;
sos_loop[0].somModel.sram_ptr[7][180]=3;
sos_loop[0].somModel.sram_dat[7][181][0]=96'h4045;
sos_loop[0].somModel.sram_ptr[7][181]=3;
sos_loop[0].somModel.sram_dat[7][182][0]=96'h2e4b;
sos_loop[0].somModel.sram_ptr[7][182]=3;
sos_loop[0].somModel.sram_dat[7][183][0]=96'h5001;
sos_loop[0].somModel.sram_ptr[7][183]=3;
sos_loop[0].somModel.sram_dat[7][184][0]=96'h89f4;
sos_loop[0].somModel.sram_ptr[7][184]=3;
sos_loop[0].somModel.sram_dat[7][185][0]=96'h4f20;
sos_loop[0].somModel.sram_ptr[7][185]=3;
sos_loop[0].somModel.sram_dat[7][186][0]=96'h718d;
sos_loop[0].somModel.sram_ptr[7][186]=3;
sos_loop[0].somModel.sram_dat[7][187][0]=96'hec81;
sos_loop[0].somModel.sram_ptr[7][187]=3;
sos_loop[0].somModel.sram_dat[7][188][0]=96'heff2;
sos_loop[0].somModel.sram_ptr[7][188]=3;
sos_loop[0].somModel.sram_dat[7][189][0]=96'h32f9;
sos_loop[0].somModel.sram_ptr[7][189]=3;
sos_loop[0].somModel.sram_dat[7][190][0]=96'hdf51;
sos_loop[0].somModel.sram_ptr[7][190]=3;
sos_loop[0].somModel.sram_dat[7][191][0]=96'haebe;
sos_loop[0].somModel.sram_ptr[7][191]=3;
sos_loop[0].somModel.sram_dat[7][192][0]=96'h1952;
sos_loop[0].somModel.sram_ptr[7][192]=3;
sos_loop[0].somModel.sram_dat[7][193][0]=96'h989a;
sos_loop[0].somModel.sram_ptr[7][193]=3;
sos_loop[0].somModel.sram_dat[7][194][0]=96'h4d90;
sos_loop[0].somModel.sram_ptr[7][194]=3;
sos_loop[0].somModel.sram_dat[7][195][0]=96'hcda6;
sos_loop[0].somModel.sram_ptr[7][195]=3;
sos_loop[0].somModel.sram_dat[7][196][0]=96'h11cf;
sos_loop[0].somModel.sram_ptr[7][196]=3;
sos_loop[0].somModel.sram_dat[7][197][0]=96'h46d5;
sos_loop[0].somModel.sram_ptr[7][197]=3;
sos_loop[0].somModel.sram_dat[7][198][0]=96'hcdeb;
sos_loop[0].somModel.sram_ptr[7][198]=3;
sos_loop[0].somModel.sram_dat[7][199][0]=96'h60b3;
sos_loop[0].somModel.sram_ptr[7][199]=3;
sos_loop[0].somModel.sram_dat[7][200][0]=96'he8cc;
sos_loop[0].somModel.sram_ptr[7][200]=3;
sos_loop[0].somModel.sram_dat[7][201][0]=96'h99ed;
sos_loop[0].somModel.sram_ptr[7][201]=3;
sos_loop[0].somModel.sram_dat[7][202][0]=96'hc9aa;
sos_loop[0].somModel.sram_ptr[7][202]=3;
sos_loop[0].somModel.sram_dat[7][203][0]=96'ha401;
sos_loop[0].somModel.sram_ptr[7][203]=3;
sos_loop[0].somModel.sram_dat[7][204][0]=96'ha4a0;
sos_loop[0].somModel.sram_ptr[7][204]=3;
sos_loop[0].somModel.sram_dat[7][205][0]=96'h9821;
sos_loop[0].somModel.sram_ptr[7][205]=3;
sos_loop[0].somModel.sram_dat[7][206][0]=96'he330;
sos_loop[0].somModel.sram_ptr[7][206]=3;
sos_loop[0].somModel.sram_dat[7][207][0]=96'h5327;
sos_loop[0].somModel.sram_ptr[7][207]=3;
sos_loop[0].somModel.sram_dat[7][208][0]=96'h85c;
sos_loop[0].somModel.sram_ptr[7][208]=3;
sos_loop[0].somModel.sram_dat[7][209][0]=96'hf8ea;
sos_loop[0].somModel.sram_ptr[7][209]=3;
sos_loop[0].somModel.sram_dat[7][210][0]=96'h243d;
sos_loop[0].somModel.sram_ptr[7][210]=3;
sos_loop[0].somModel.sram_dat[7][211][0]=96'h67f8;
sos_loop[0].somModel.sram_ptr[7][211]=3;
sos_loop[0].somModel.sram_dat[7][212][0]=96'h55bf;
sos_loop[0].somModel.sram_ptr[7][212]=3;
sos_loop[0].somModel.sram_dat[7][213][0]=96'h731b;
sos_loop[0].somModel.sram_ptr[7][213]=3;
sos_loop[0].somModel.sram_dat[7][214][0]=96'h80fd;
sos_loop[0].somModel.sram_ptr[7][214]=3;
sos_loop[0].somModel.sram_dat[7][215][0]=96'haf4c;
sos_loop[0].somModel.sram_ptr[7][215]=3;
sos_loop[0].somModel.sram_dat[7][216][0]=96'h4a57;
sos_loop[0].somModel.sram_ptr[7][216]=3;
sos_loop[0].somModel.sram_dat[7][217][0]=96'h414d;
sos_loop[0].somModel.sram_ptr[7][217]=3;
sos_loop[0].somModel.sram_dat[7][218][0]=96'h5dd0;
sos_loop[0].somModel.sram_ptr[7][218]=3;
sos_loop[0].somModel.sram_dat[7][219][0]=96'h7720;
sos_loop[0].somModel.sram_ptr[7][219]=3;
sos_loop[0].somModel.sram_dat[7][220][0]=96'h378c;
sos_loop[0].somModel.sram_ptr[7][220]=3;
sos_loop[0].somModel.sram_dat[7][221][0]=96'hc49c;
sos_loop[0].somModel.sram_ptr[7][221]=3;
sos_loop[0].somModel.sram_dat[7][222][0]=96'h97f4;
sos_loop[0].somModel.sram_ptr[7][222]=3;
sos_loop[0].somModel.sram_dat[7][223][0]=96'h7335;
sos_loop[0].somModel.sram_ptr[7][223]=3;
sos_loop[0].somModel.sram_dat[7][224][0]=96'h130f;
sos_loop[0].somModel.sram_ptr[7][224]=3;
sos_loop[0].somModel.sram_dat[7][225][0]=96'h9dc0;
sos_loop[0].somModel.sram_ptr[7][225]=3;
sos_loop[0].somModel.sram_dat[7][226][0]=96'hf760;
sos_loop[0].somModel.sram_ptr[7][226]=3;
sos_loop[0].somModel.sram_dat[7][227][0]=96'h1800;
sos_loop[0].somModel.sram_ptr[7][227]=3;
sos_loop[0].somModel.sram_dat[7][228][0]=96'h40fe;
sos_loop[0].somModel.sram_ptr[7][228]=3;
sos_loop[0].somModel.sram_dat[7][229][0]=96'h698d;
sos_loop[0].somModel.sram_ptr[7][229]=3;
sos_loop[0].somModel.sram_dat[7][230][0]=96'hac63;
sos_loop[0].somModel.sram_ptr[7][230]=3;
sos_loop[0].somModel.sram_dat[7][231][0]=96'hcb0;
sos_loop[0].somModel.sram_ptr[7][231]=3;
sos_loop[0].somModel.sram_dat[7][232][0]=96'ha762;
sos_loop[0].somModel.sram_ptr[7][232]=3;
sos_loop[0].somModel.sram_dat[7][233][0]=96'hc7e3;
sos_loop[0].somModel.sram_ptr[7][233]=3;
sos_loop[0].somModel.sram_dat[7][234][0]=96'h7950;
sos_loop[0].somModel.sram_ptr[7][234]=3;
sos_loop[0].somModel.sram_dat[7][235][0]=96'h393f;
sos_loop[0].somModel.sram_ptr[7][235]=3;
sos_loop[0].somModel.sram_dat[7][236][0]=96'hb5a0;
sos_loop[0].somModel.sram_ptr[7][236]=3;
sos_loop[0].somModel.sram_dat[7][237][0]=96'ha992;
sos_loop[0].somModel.sram_ptr[7][237]=3;
sos_loop[0].somModel.sram_dat[7][238][0]=96'h9d82;
sos_loop[0].somModel.sram_ptr[7][238]=3;
sos_loop[0].somModel.sram_dat[7][239][0]=96'h4659;
sos_loop[0].somModel.sram_ptr[7][239]=3;
sos_loop[0].somModel.sram_dat[7][240][0]=96'h99f3;
sos_loop[0].somModel.sram_ptr[7][240]=3;
sos_loop[0].somModel.sram_dat[7][241][0]=96'h31f6;
sos_loop[0].somModel.sram_ptr[7][241]=3;
sos_loop[0].somModel.sram_dat[7][242][0]=96'h4389;
sos_loop[0].somModel.sram_ptr[7][242]=3;
sos_loop[0].somModel.sram_dat[7][243][0]=96'h9fbe;
sos_loop[0].somModel.sram_ptr[7][243]=3;
sos_loop[0].somModel.sram_dat[7][244][0]=96'h1fa1;
sos_loop[0].somModel.sram_ptr[7][244]=3;
sos_loop[0].somModel.sram_dat[7][245][0]=96'h4eb0;
sos_loop[0].somModel.sram_ptr[7][245]=3;
sos_loop[0].somModel.sram_dat[7][246][0]=96'haf41;
sos_loop[0].somModel.sram_ptr[7][246]=3;
sos_loop[0].somModel.sram_dat[7][247][0]=96'h8b0d;
sos_loop[0].somModel.sram_ptr[7][247]=3;
sos_loop[0].somModel.sram_dat[7][248][0]=96'hb721;
sos_loop[0].somModel.sram_ptr[7][248]=3;
sos_loop[0].somModel.sram_dat[7][249][0]=96'hb055;
sos_loop[0].somModel.sram_ptr[7][249]=3;
sos_loop[0].somModel.sram_dat[7][250][0]=96'ha3fa;
sos_loop[0].somModel.sram_ptr[7][250]=3;
sos_loop[0].somModel.sram_dat[7][251][0]=96'hf530;
sos_loop[0].somModel.sram_ptr[7][251]=3;
sos_loop[0].somModel.sram_dat[7][252][0]=96'h40ec;
sos_loop[0].somModel.sram_ptr[7][252]=3;
sos_loop[0].somModel.sram_dat[7][253][0]=96'hbf82;
sos_loop[0].somModel.sram_ptr[7][253]=3;
sos_loop[0].somModel.sram_dat[7][254][0]=96'h2613;
sos_loop[0].somModel.sram_ptr[7][254]=3;
sos_loop[0].somModel.sram_dat[7][255][0]=96'h7010;
sos_loop[0].somModel.sram_ptr[7][255]=3;
sos_loop[0].somModel.sram_dat[7][256][0]=96'hc20c;
sos_loop[0].somModel.sram_ptr[7][256]=3;
sos_loop[0].somModel.sram_dat[7][257][0]=96'hb5a2;
sos_loop[0].somModel.sram_ptr[7][257]=3;
sos_loop[0].somModel.sram_dat[7][258][0]=96'h7d6;
sos_loop[0].somModel.sram_ptr[7][258]=3;
sos_loop[0].somModel.sram_dat[7][259][0]=96'h8c9b;
sos_loop[0].somModel.sram_ptr[7][259]=3;
sos_loop[0].somModel.sram_dat[7][260][0]=96'h2cb2;
sos_loop[0].somModel.sram_ptr[7][260]=3;
sos_loop[0].somModel.sram_dat[7][261][0]=96'hac1b;
sos_loop[0].somModel.sram_ptr[7][261]=3;
sos_loop[0].somModel.sram_dat[7][262][0]=96'hc493;
sos_loop[0].somModel.sram_ptr[7][262]=3;
sos_loop[0].somModel.sram_dat[7][263][0]=96'h2fc6;
sos_loop[0].somModel.sram_ptr[7][263]=3;
sos_loop[0].somModel.sram_dat[7][264][0]=96'ha2b9;
sos_loop[0].somModel.sram_ptr[7][264]=3;
sos_loop[0].somModel.sram_dat[7][265][0]=96'hf03a;
sos_loop[0].somModel.sram_ptr[7][265]=3;
sos_loop[0].somModel.sram_dat[7][266][0]=96'h628c;
sos_loop[0].somModel.sram_ptr[7][266]=3;
sos_loop[0].somModel.sram_dat[7][267][0]=96'h8a4f;
sos_loop[0].somModel.sram_ptr[7][267]=3;
sos_loop[0].somModel.sram_dat[7][268][0]=96'hf6ce;
sos_loop[0].somModel.sram_ptr[7][268]=3;
sos_loop[0].somModel.sram_dat[7][269][0]=96'h94f6;
sos_loop[0].somModel.sram_ptr[7][269]=3;
sos_loop[0].somModel.sram_dat[7][270][0]=96'h5ff0;
sos_loop[0].somModel.sram_ptr[7][270]=3;
sos_loop[0].somModel.sram_dat[7][271][0]=96'hdd7f;
sos_loop[0].somModel.sram_ptr[7][271]=3;
sos_loop[0].somModel.sram_dat[7][272][0]=96'he12f;
sos_loop[0].somModel.sram_ptr[7][272]=3;
sos_loop[0].somModel.sram_dat[7][273][0]=96'h773e;
sos_loop[0].somModel.sram_ptr[7][273]=3;
sos_loop[0].somModel.sram_dat[7][274][0]=96'hadd4;
sos_loop[0].somModel.sram_ptr[7][274]=3;
sos_loop[0].somModel.sram_dat[7][275][0]=96'hbc61;
sos_loop[0].somModel.sram_ptr[7][275]=3;
sos_loop[0].somModel.sram_dat[7][276][0]=96'hbce1;
sos_loop[0].somModel.sram_ptr[7][276]=3;
sos_loop[0].somModel.sram_dat[7][277][0]=96'h7c3d;
sos_loop[0].somModel.sram_ptr[7][277]=3;
sos_loop[0].somModel.sram_dat[7][278][0]=96'hcbb3;
sos_loop[0].somModel.sram_ptr[7][278]=3;
sos_loop[0].somModel.sram_dat[7][279][0]=96'h47e1;
sos_loop[0].somModel.sram_ptr[7][279]=3;
sos_loop[0].somModel.sram_dat[7][280][0]=96'h54ac;
sos_loop[0].somModel.sram_ptr[7][280]=3;
sos_loop[0].somModel.sram_dat[7][281][0]=96'hd99;
sos_loop[0].somModel.sram_ptr[7][281]=3;
sos_loop[0].somModel.sram_dat[7][282][0]=96'h337c;
sos_loop[0].somModel.sram_ptr[7][282]=3;
sos_loop[0].somModel.sram_dat[7][283][0]=96'h70b8;
sos_loop[0].somModel.sram_ptr[7][283]=3;
sos_loop[0].somModel.sram_dat[7][284][0]=96'h732e;
sos_loop[0].somModel.sram_ptr[7][284]=3;
sos_loop[0].somModel.sram_dat[7][285][0]=96'h6d44;
sos_loop[0].somModel.sram_ptr[7][285]=3;
sos_loop[0].somModel.sram_dat[7][286][0]=96'h5f66;
sos_loop[0].somModel.sram_ptr[7][286]=3;
sos_loop[0].somModel.sram_dat[7][287][0]=96'hcead;
sos_loop[0].somModel.sram_ptr[7][287]=3;
sos_loop[0].somModel.sram_dat[7][288][0]=96'h35a7;
sos_loop[0].somModel.sram_ptr[7][288]=3;
sos_loop[0].somModel.sram_dat[7][289][0]=96'h36bd;
sos_loop[0].somModel.sram_ptr[7][289]=3;
sos_loop[0].somModel.sram_dat[7][290][0]=96'h9924;
sos_loop[0].somModel.sram_ptr[7][290]=3;
sos_loop[0].somModel.sram_dat[7][291][0]=96'h9e17;
sos_loop[0].somModel.sram_ptr[7][291]=3;
sos_loop[0].somModel.sram_dat[7][292][0]=96'hc72a;
sos_loop[0].somModel.sram_ptr[7][292]=3;
sos_loop[0].somModel.sram_dat[7][293][0]=96'h4ee3;
sos_loop[0].somModel.sram_ptr[7][293]=3;
sos_loop[0].somModel.sram_dat[7][294][0]=96'h5e7;
sos_loop[0].somModel.sram_ptr[7][294]=3;
sos_loop[0].somModel.sram_dat[7][295][0]=96'hb1e7;
sos_loop[0].somModel.sram_ptr[7][295]=3;
sos_loop[0].somModel.sram_dat[7][296][0]=96'h5cac;
sos_loop[0].somModel.sram_ptr[7][296]=3;
sos_loop[0].somModel.sram_dat[7][297][0]=96'h7c98;
sos_loop[0].somModel.sram_ptr[7][297]=3;
sos_loop[0].somModel.sram_dat[7][298][0]=96'hf24a;
sos_loop[0].somModel.sram_ptr[7][298]=3;
sos_loop[0].somModel.sram_dat[7][299][0]=96'h9017;
sos_loop[0].somModel.sram_ptr[7][299]=3;
sos_loop[0].somModel.sram_dat[7][300][0]=96'ha86;
sos_loop[0].somModel.sram_ptr[7][300]=3;
sos_loop[0].somModel.sram_dat[7][301][0]=96'h15c7;
sos_loop[0].somModel.sram_ptr[7][301]=3;
sos_loop[0].somModel.sram_dat[7][302][0]=96'h6c3d;
sos_loop[0].somModel.sram_ptr[7][302]=3;
sos_loop[0].somModel.sram_dat[7][303][0]=96'h501e;
sos_loop[0].somModel.sram_ptr[7][303]=3;
sos_loop[0].somModel.sram_dat[7][304][0]=96'h10c9;
sos_loop[0].somModel.sram_ptr[7][304]=3;
sos_loop[0].somModel.sram_dat[7][305][0]=96'h5862;
sos_loop[0].somModel.sram_ptr[7][305]=3;
sos_loop[0].somModel.sram_dat[7][306][0]=96'h28e;
sos_loop[0].somModel.sram_ptr[7][306]=3;
sos_loop[0].somModel.sram_dat[7][307][0]=96'hc850;
sos_loop[0].somModel.sram_ptr[7][307]=3;
sos_loop[0].somModel.sram_dat[7][308][0]=96'haf6c;
sos_loop[0].somModel.sram_ptr[7][308]=3;
sos_loop[0].somModel.sram_dat[7][309][0]=96'h90d3;
sos_loop[0].somModel.sram_ptr[7][309]=3;
sos_loop[0].somModel.sram_dat[7][310][0]=96'hb6b1;
sos_loop[0].somModel.sram_ptr[7][310]=3;
sos_loop[0].somModel.sram_dat[7][311][0]=96'h5e8d;
sos_loop[0].somModel.sram_ptr[7][311]=3;
sos_loop[0].somModel.sram_dat[7][312][0]=96'h5855;
sos_loop[0].somModel.sram_ptr[7][312]=3;
sos_loop[0].somModel.sram_dat[7][313][0]=96'h6c01;
sos_loop[0].somModel.sram_ptr[7][313]=3;
sos_loop[0].somModel.sram_dat[7][314][0]=96'hdcb4;
sos_loop[0].somModel.sram_ptr[7][314]=3;
sos_loop[0].somModel.sram_dat[7][315][0]=96'hc207;
sos_loop[0].somModel.sram_ptr[7][315]=3;
sos_loop[0].somModel.sram_dat[7][316][0]=96'hf4c7;
sos_loop[0].somModel.sram_ptr[7][316]=3;
sos_loop[0].somModel.sram_dat[7][317][0]=96'hc655;
sos_loop[0].somModel.sram_ptr[7][317]=3;
sos_loop[0].somModel.sram_dat[7][318][0]=96'h5a6a;
sos_loop[0].somModel.sram_ptr[7][318]=3;
sos_loop[0].somModel.sram_dat[7][319][0]=96'hfdf1;
sos_loop[0].somModel.sram_ptr[7][319]=3;
sos_loop[0].somModel.sram_dat[7][320][0]=96'h762c;
sos_loop[0].somModel.sram_ptr[7][320]=3;
sos_loop[0].somModel.sram_dat[7][321][0]=96'h3342;
sos_loop[0].somModel.sram_ptr[7][321]=3;
sos_loop[0].somModel.sram_dat[7][322][0]=96'ha47d;
sos_loop[0].somModel.sram_ptr[7][322]=3;
sos_loop[0].somModel.sram_dat[7][323][0]=96'h49d;
sos_loop[0].somModel.sram_ptr[7][323]=3;
sos_loop[0].somModel.sram_dat[7][324][0]=96'h4c88;
sos_loop[0].somModel.sram_ptr[7][324]=3;
sos_loop[0].somModel.sram_dat[7][325][0]=96'hb9a2;
sos_loop[0].somModel.sram_ptr[7][325]=3;
sos_loop[0].somModel.sram_dat[7][326][0]=96'h605b;
sos_loop[0].somModel.sram_ptr[7][326]=3;
sos_loop[0].somModel.sram_dat[7][327][0]=96'h1b57;
sos_loop[0].somModel.sram_ptr[7][327]=3;
sos_loop[0].somModel.sram_dat[7][328][0]=96'h2d7c;
sos_loop[0].somModel.sram_ptr[7][328]=3;
sos_loop[0].somModel.sram_dat[7][329][0]=96'h598d;
sos_loop[0].somModel.sram_ptr[7][329]=3;
sos_loop[0].somModel.sram_dat[7][330][0]=96'hbad0;
sos_loop[0].somModel.sram_ptr[7][330]=3;
sos_loop[0].somModel.sram_dat[7][331][0]=96'h2246;
sos_loop[0].somModel.sram_ptr[7][331]=3;
sos_loop[0].somModel.sram_dat[7][332][0]=96'ha559;
sos_loop[0].somModel.sram_ptr[7][332]=3;
sos_loop[0].somModel.sram_dat[7][333][0]=96'he9bd;
sos_loop[0].somModel.sram_ptr[7][333]=3;
sos_loop[0].somModel.sram_dat[7][334][0]=96'hba7c;
sos_loop[0].somModel.sram_ptr[7][334]=3;
sos_loop[0].somModel.sram_dat[7][335][0]=96'hbf4e;
sos_loop[0].somModel.sram_ptr[7][335]=3;
sos_loop[0].somModel.sram_dat[7][336][0]=96'h505a;
sos_loop[0].somModel.sram_ptr[7][336]=3;
sos_loop[0].somModel.sram_dat[7][337][0]=96'h7213;
sos_loop[0].somModel.sram_ptr[7][337]=3;
sos_loop[0].somModel.sram_dat[7][338][0]=96'h7e6d;
sos_loop[0].somModel.sram_ptr[7][338]=3;
sos_loop[0].somModel.sram_dat[7][339][0]=96'h676e;
sos_loop[0].somModel.sram_ptr[7][339]=3;
sos_loop[0].somModel.sram_dat[7][340][0]=96'h191f;
sos_loop[0].somModel.sram_ptr[7][340]=3;
sos_loop[0].somModel.sram_dat[7][341][0]=96'h3181;
sos_loop[0].somModel.sram_ptr[7][341]=3;
sos_loop[0].somModel.sram_dat[7][342][0]=96'h17ab;
sos_loop[0].somModel.sram_ptr[7][342]=3;
sos_loop[0].somModel.sram_dat[7][343][0]=96'h3075;
sos_loop[0].somModel.sram_ptr[7][343]=3;
sos_loop[0].somModel.sram_dat[7][344][0]=96'hafc7;
sos_loop[0].somModel.sram_ptr[7][344]=3;
sos_loop[0].somModel.sram_dat[7][345][0]=96'hcde1;
sos_loop[0].somModel.sram_ptr[7][345]=3;
sos_loop[0].somModel.sram_dat[7][346][0]=96'h4ffc;
sos_loop[0].somModel.sram_ptr[7][346]=3;
sos_loop[0].somModel.sram_dat[7][347][0]=96'hdc23;
sos_loop[0].somModel.sram_ptr[7][347]=3;
sos_loop[0].somModel.sram_dat[7][348][0]=96'hd21;
sos_loop[0].somModel.sram_ptr[7][348]=3;
sos_loop[0].somModel.sram_dat[7][349][0]=96'h6432;
sos_loop[0].somModel.sram_ptr[7][349]=3;
sos_loop[0].somModel.sram_dat[7][350][0]=96'h925a;
sos_loop[0].somModel.sram_ptr[7][350]=3;
sos_loop[0].somModel.sram_dat[7][351][0]=96'hc72e;
sos_loop[0].somModel.sram_ptr[7][351]=3;
sos_loop[0].somModel.sram_dat[7][352][0]=96'h59d9;
sos_loop[0].somModel.sram_ptr[7][352]=3;
sos_loop[0].somModel.sram_dat[7][353][0]=96'h7e41;
sos_loop[0].somModel.sram_ptr[7][353]=3;
sos_loop[0].somModel.sram_dat[7][354][0]=96'he51e;
sos_loop[0].somModel.sram_ptr[7][354]=3;
sos_loop[0].somModel.sram_dat[7][355][0]=96'h2182;
sos_loop[0].somModel.sram_ptr[7][355]=3;
sos_loop[0].somModel.sram_dat[7][356][0]=96'h85fd;
sos_loop[0].somModel.sram_ptr[7][356]=3;
sos_loop[0].somModel.sram_dat[7][357][0]=96'hff81;
sos_loop[0].somModel.sram_ptr[7][357]=3;
sos_loop[0].somModel.sram_dat[7][358][0]=96'habc8;
sos_loop[0].somModel.sram_ptr[7][358]=3;
sos_loop[0].somModel.sram_dat[7][359][0]=96'h933;
sos_loop[0].somModel.sram_ptr[7][359]=3;
sos_loop[0].somModel.sram_dat[7][360][0]=96'h75b;
sos_loop[0].somModel.sram_ptr[7][360]=3;
sos_loop[0].somModel.sram_dat[7][361][0]=96'he194;
sos_loop[0].somModel.sram_ptr[7][361]=3;
sos_loop[0].somModel.sram_dat[7][362][0]=96'ha000;
sos_loop[0].somModel.sram_ptr[7][362]=3;
sos_loop[0].somModel.sram_dat[7][363][0]=96'h75d7;
sos_loop[0].somModel.sram_ptr[7][363]=3;
sos_loop[0].somModel.sram_dat[7][364][0]=96'h2796;
sos_loop[0].somModel.sram_ptr[7][364]=3;
sos_loop[0].somModel.sram_dat[7][365][0]=96'he2de;
sos_loop[0].somModel.sram_ptr[7][365]=3;
sos_loop[0].somModel.sram_dat[7][366][0]=96'hfb48;
sos_loop[0].somModel.sram_ptr[7][366]=3;
sos_loop[0].somModel.sram_dat[7][367][0]=96'h6be4;
sos_loop[0].somModel.sram_ptr[7][367]=3;
sos_loop[0].somModel.sram_dat[7][368][0]=96'ha2f;
sos_loop[0].somModel.sram_ptr[7][368]=3;
sos_loop[0].somModel.sram_dat[7][369][0]=96'h8b4f;
sos_loop[0].somModel.sram_ptr[7][369]=3;
sos_loop[0].somModel.sram_dat[7][370][0]=96'hf592;
sos_loop[0].somModel.sram_ptr[7][370]=3;
sos_loop[0].somModel.sram_dat[7][371][0]=96'h2cc7;
sos_loop[0].somModel.sram_ptr[7][371]=3;
sos_loop[0].somModel.sram_dat[7][372][0]=96'hb053;
sos_loop[0].somModel.sram_ptr[7][372]=3;
sos_loop[0].somModel.sram_dat[7][373][0]=96'ha982;
sos_loop[0].somModel.sram_ptr[7][373]=3;
sos_loop[0].somModel.sram_dat[7][374][0]=96'hf7f5;
sos_loop[0].somModel.sram_ptr[7][374]=3;
sos_loop[0].somModel.sram_dat[7][375][0]=96'habff;
sos_loop[0].somModel.sram_ptr[7][375]=3;
sos_loop[0].somModel.sram_dat[7][376][0]=96'hc5a1;
sos_loop[0].somModel.sram_ptr[7][376]=3;
sos_loop[0].somModel.sram_dat[7][377][0]=96'hc504;
sos_loop[0].somModel.sram_ptr[7][377]=3;
sos_loop[0].somModel.sram_dat[7][378][0]=96'h260b;
sos_loop[0].somModel.sram_ptr[7][378]=3;
sos_loop[0].somModel.sram_dat[7][379][0]=96'hecef;
sos_loop[0].somModel.sram_ptr[7][379]=3;
sos_loop[0].somModel.sram_dat[7][380][0]=96'h1548;
sos_loop[0].somModel.sram_ptr[7][380]=3;
sos_loop[0].somModel.sram_dat[7][381][0]=96'h63f7;
sos_loop[0].somModel.sram_ptr[7][381]=3;
sos_loop[0].somModel.sram_dat[7][382][0]=96'h97c;
sos_loop[0].somModel.sram_ptr[7][382]=3;
sos_loop[0].somModel.sram_dat[7][383][0]=96'h492e;
sos_loop[0].somModel.sram_ptr[7][383]=3;
sos_loop[0].somModel.sram_dat[7][384][0]=96'h7d91;
sos_loop[0].somModel.sram_ptr[7][384]=3;
sos_loop[0].somModel.sram_dat[7][385][0]=96'h5e33;
sos_loop[0].somModel.sram_ptr[7][385]=3;
sos_loop[0].somModel.sram_dat[7][386][0]=96'h20ff;
sos_loop[0].somModel.sram_ptr[7][386]=3;
sos_loop[0].somModel.sram_dat[7][387][0]=96'h2d2b;
sos_loop[0].somModel.sram_ptr[7][387]=3;
sos_loop[0].somModel.sram_dat[7][388][0]=96'h4faf;
sos_loop[0].somModel.sram_ptr[7][388]=3;
sos_loop[0].somModel.sram_dat[7][389][0]=96'h9fc0;
sos_loop[0].somModel.sram_ptr[7][389]=3;
sos_loop[0].somModel.sram_dat[7][390][0]=96'h7df6;
sos_loop[0].somModel.sram_ptr[7][390]=3;
sos_loop[0].somModel.sram_dat[7][391][0]=96'h8145;
sos_loop[0].somModel.sram_ptr[7][391]=3;
sos_loop[0].somModel.sram_dat[7][392][0]=96'hd8dc;
sos_loop[0].somModel.sram_ptr[7][392]=3;
sos_loop[0].somModel.sram_dat[7][393][0]=96'h8ccb;
sos_loop[0].somModel.sram_ptr[7][393]=3;
sos_loop[0].somModel.sram_dat[7][394][0]=96'ha74c;
sos_loop[0].somModel.sram_ptr[7][394]=3;
sos_loop[0].somModel.sram_dat[7][395][0]=96'hd54d;
sos_loop[0].somModel.sram_ptr[7][395]=3;
sos_loop[0].somModel.sram_dat[7][396][0]=96'h57ec;
sos_loop[0].somModel.sram_ptr[7][396]=3;
sos_loop[0].somModel.sram_dat[7][397][0]=96'hd895;
sos_loop[0].somModel.sram_ptr[7][397]=3;
sos_loop[0].somModel.sram_dat[7][398][0]=96'h4a8a;
sos_loop[0].somModel.sram_ptr[7][398]=3;
sos_loop[0].somModel.sram_dat[7][399][0]=96'haad5;
sos_loop[0].somModel.sram_ptr[7][399]=3;
sos_loop[0].somModel.sram_dat[7][400][0]=96'h2dc8;
sos_loop[0].somModel.sram_ptr[7][400]=3;
sos_loop[0].somModel.sram_dat[7][401][0]=96'hd305;
sos_loop[0].somModel.sram_ptr[7][401]=3;
sos_loop[0].somModel.sram_dat[7][402][0]=96'hf654;
sos_loop[0].somModel.sram_ptr[7][402]=3;
sos_loop[0].somModel.sram_dat[7][403][0]=96'h7cef;
sos_loop[0].somModel.sram_ptr[7][403]=3;
sos_loop[0].somModel.sram_dat[7][404][0]=96'hfdcd;
sos_loop[0].somModel.sram_ptr[7][404]=3;
sos_loop[0].somModel.sram_dat[7][405][0]=96'h9c53;
sos_loop[0].somModel.sram_ptr[7][405]=3;
sos_loop[0].somModel.sram_dat[7][406][0]=96'h56bf;
sos_loop[0].somModel.sram_ptr[7][406]=3;
sos_loop[0].somModel.sram_dat[7][407][0]=96'hdf03;
sos_loop[0].somModel.sram_ptr[7][407]=3;
sos_loop[0].somModel.sram_dat[7][408][0]=96'h8eb7;
sos_loop[0].somModel.sram_ptr[7][408]=3;
sos_loop[0].somModel.sram_dat[7][409][0]=96'h27c4;
sos_loop[0].somModel.sram_ptr[7][409]=3;
sos_loop[0].somModel.sram_dat[7][410][0]=96'h6ae4;
sos_loop[0].somModel.sram_ptr[7][410]=3;
sos_loop[0].somModel.sram_dat[7][411][0]=96'h8beb;
sos_loop[0].somModel.sram_ptr[7][411]=3;
sos_loop[0].somModel.sram_dat[7][412][0]=96'h6ac7;
sos_loop[0].somModel.sram_ptr[7][412]=3;
sos_loop[0].somModel.sram_dat[7][413][0]=96'hc8ce;
sos_loop[0].somModel.sram_ptr[7][413]=3;
sos_loop[0].somModel.sram_dat[7][414][0]=96'hf6f;
sos_loop[0].somModel.sram_ptr[7][414]=3;
sos_loop[0].somModel.sram_dat[7][415][0]=96'hc185;
sos_loop[0].somModel.sram_ptr[7][415]=3;
sos_loop[0].somModel.sram_dat[7][416][0]=96'h8ecb;
sos_loop[0].somModel.sram_ptr[7][416]=3;
sos_loop[0].somModel.sram_dat[7][417][0]=96'hc088;
sos_loop[0].somModel.sram_ptr[7][417]=3;
sos_loop[0].somModel.sram_dat[7][418][0]=96'hfb13;
sos_loop[0].somModel.sram_ptr[7][418]=3;
sos_loop[0].somModel.sram_dat[7][419][0]=96'h8323;
sos_loop[0].somModel.sram_ptr[7][419]=3;
sos_loop[0].somModel.sram_dat[7][420][0]=96'h4be;
sos_loop[0].somModel.sram_ptr[7][420]=3;
sos_loop[0].somModel.sram_dat[7][421][0]=96'hd5d8;
sos_loop[0].somModel.sram_ptr[7][421]=3;
sos_loop[0].somModel.sram_dat[7][422][0]=96'hf5e5;
sos_loop[0].somModel.sram_ptr[7][422]=3;
sos_loop[0].somModel.sram_dat[7][423][0]=96'he858;
sos_loop[0].somModel.sram_ptr[7][423]=3;
sos_loop[0].somModel.sram_dat[7][424][0]=96'hec83;
sos_loop[0].somModel.sram_ptr[7][424]=3;
sos_loop[0].somModel.sram_dat[7][425][0]=96'h4b57;
sos_loop[0].somModel.sram_ptr[7][425]=3;
sos_loop[0].somModel.sram_dat[7][426][0]=96'h7510;
sos_loop[0].somModel.sram_ptr[7][426]=3;
sos_loop[0].somModel.sram_dat[7][427][0]=96'h7e0c;
sos_loop[0].somModel.sram_ptr[7][427]=3;
sos_loop[0].somModel.sram_dat[7][428][0]=96'hafdd;
sos_loop[0].somModel.sram_ptr[7][428]=3;
sos_loop[0].somModel.sram_dat[7][429][0]=96'heea0;
sos_loop[0].somModel.sram_ptr[7][429]=3;
sos_loop[0].somModel.sram_dat[7][430][0]=96'hdc6b;
sos_loop[0].somModel.sram_ptr[7][430]=3;
sos_loop[0].somModel.sram_dat[7][431][0]=96'hdc6d;
sos_loop[0].somModel.sram_ptr[7][431]=3;
sos_loop[0].somModel.sram_dat[7][432][0]=96'hf267;
sos_loop[0].somModel.sram_ptr[7][432]=3;
sos_loop[0].somModel.sram_dat[7][433][0]=96'hcc96;
sos_loop[0].somModel.sram_ptr[7][433]=3;
sos_loop[0].somModel.sram_dat[7][434][0]=96'h6e0e;
sos_loop[0].somModel.sram_ptr[7][434]=3;
sos_loop[0].somModel.sram_dat[7][435][0]=96'hadf2;
sos_loop[0].somModel.sram_ptr[7][435]=3;
sos_loop[0].somModel.sram_dat[7][436][0]=96'h22cf;
sos_loop[0].somModel.sram_ptr[7][436]=3;
sos_loop[0].somModel.sram_dat[7][437][0]=96'hefe3;
sos_loop[0].somModel.sram_ptr[7][437]=3;
sos_loop[0].somModel.sram_dat[7][438][0]=96'h327f;
sos_loop[0].somModel.sram_ptr[7][438]=3;
sos_loop[0].somModel.sram_dat[7][439][0]=96'hc1cd;
sos_loop[0].somModel.sram_ptr[7][439]=3;
sos_loop[0].somModel.sram_dat[7][440][0]=96'h87d7;
sos_loop[0].somModel.sram_ptr[7][440]=3;
sos_loop[0].somModel.sram_dat[7][441][0]=96'h52ae;
sos_loop[0].somModel.sram_ptr[7][441]=3;
sos_loop[0].somModel.sram_dat[7][442][0]=96'h522d;
sos_loop[0].somModel.sram_ptr[7][442]=3;
sos_loop[0].somModel.sram_dat[7][443][0]=96'h23e9;
sos_loop[0].somModel.sram_ptr[7][443]=3;
sos_loop[0].somModel.sram_dat[7][444][0]=96'h9f00;
sos_loop[0].somModel.sram_ptr[7][444]=3;
sos_loop[0].somModel.sram_dat[7][445][0]=96'h4222;
sos_loop[0].somModel.sram_ptr[7][445]=3;
sos_loop[0].somModel.sram_dat[7][446][0]=96'hc826;
sos_loop[0].somModel.sram_ptr[7][446]=3;
sos_loop[0].somModel.sram_dat[7][447][0]=96'h5c33;
sos_loop[0].somModel.sram_ptr[7][447]=3;
sos_loop[0].somModel.sram_dat[7][448][0]=96'h25c2;
sos_loop[0].somModel.sram_ptr[7][448]=3;
sos_loop[0].somModel.sram_dat[7][449][0]=96'hc4f6;
sos_loop[0].somModel.sram_ptr[7][449]=3;
sos_loop[0].somModel.sram_dat[7][450][0]=96'hf947;
sos_loop[0].somModel.sram_ptr[7][450]=3;
sos_loop[0].somModel.sram_dat[7][451][0]=96'h75e1;
sos_loop[0].somModel.sram_ptr[7][451]=3;
sos_loop[0].somModel.sram_dat[7][452][0]=96'h4b59;
sos_loop[0].somModel.sram_ptr[7][452]=3;
sos_loop[0].somModel.sram_dat[7][453][0]=96'hcc5d;
sos_loop[0].somModel.sram_ptr[7][453]=3;
sos_loop[0].somModel.sram_dat[7][454][0]=96'hec89;
sos_loop[0].somModel.sram_ptr[7][454]=3;
sos_loop[0].somModel.sram_dat[7][455][0]=96'hac8e;
sos_loop[0].somModel.sram_ptr[7][455]=3;
sos_loop[0].somModel.sram_dat[7][456][0]=96'h9306;
sos_loop[0].somModel.sram_ptr[7][456]=3;
sos_loop[0].somModel.sram_dat[7][457][0]=96'hb015;
sos_loop[0].somModel.sram_ptr[7][457]=3;
sos_loop[0].somModel.sram_dat[7][458][0]=96'h9893;
sos_loop[0].somModel.sram_ptr[7][458]=3;
sos_loop[0].somModel.sram_dat[7][459][0]=96'ha323;
sos_loop[0].somModel.sram_ptr[7][459]=3;
sos_loop[0].somModel.sram_dat[7][460][0]=96'h2482;
sos_loop[0].somModel.sram_ptr[7][460]=3;
sos_loop[0].somModel.sram_dat[7][461][0]=96'h73ba;
sos_loop[0].somModel.sram_ptr[7][461]=3;
sos_loop[0].somModel.sram_dat[7][462][0]=96'h8241;
sos_loop[0].somModel.sram_ptr[7][462]=3;
sos_loop[0].somModel.sram_dat[7][463][0]=96'h2c7;
sos_loop[0].somModel.sram_ptr[7][463]=3;
sos_loop[0].somModel.sram_dat[7][464][0]=96'h3d42;
sos_loop[0].somModel.sram_ptr[7][464]=3;
sos_loop[0].somModel.sram_dat[7][465][0]=96'h9b8;
sos_loop[0].somModel.sram_ptr[7][465]=3;
sos_loop[0].somModel.sram_dat[7][466][0]=96'h6583;
sos_loop[0].somModel.sram_ptr[7][466]=3;
sos_loop[0].somModel.sram_dat[7][467][0]=96'he989;
sos_loop[0].somModel.sram_ptr[7][467]=3;
sos_loop[0].somModel.sram_dat[7][468][0]=96'h77b8;
sos_loop[0].somModel.sram_ptr[7][468]=3;
sos_loop[0].somModel.sram_dat[7][469][0]=96'h372f;
sos_loop[0].somModel.sram_ptr[7][469]=3;
sos_loop[0].somModel.sram_dat[7][470][0]=96'hef75;
sos_loop[0].somModel.sram_ptr[7][470]=3;
sos_loop[0].somModel.sram_dat[7][471][0]=96'he2a0;
sos_loop[0].somModel.sram_ptr[7][471]=3;
sos_loop[0].somModel.sram_dat[7][472][0]=96'hf84a;
sos_loop[0].somModel.sram_ptr[7][472]=3;
sos_loop[0].somModel.sram_dat[7][473][0]=96'he2f5;
sos_loop[0].somModel.sram_ptr[7][473]=3;
sos_loop[0].somModel.sram_dat[7][474][0]=96'hca43;
sos_loop[0].somModel.sram_ptr[7][474]=3;
sos_loop[0].somModel.sram_dat[7][475][0]=96'hb85f;
sos_loop[0].somModel.sram_ptr[7][475]=3;
sos_loop[0].somModel.sram_dat[7][476][0]=96'hb9fd;
sos_loop[0].somModel.sram_ptr[7][476]=3;
sos_loop[0].somModel.sram_dat[7][477][0]=96'h730d;
sos_loop[0].somModel.sram_ptr[7][477]=3;
sos_loop[0].somModel.sram_dat[7][478][0]=96'hbd98;
sos_loop[0].somModel.sram_ptr[7][478]=3;
sos_loop[0].somModel.sram_dat[7][479][0]=96'h7046;
sos_loop[0].somModel.sram_ptr[7][479]=3;
sos_loop[0].somModel.sram_dat[7][480][0]=96'hc7f0;
sos_loop[0].somModel.sram_ptr[7][480]=3;
sos_loop[0].somModel.sram_dat[7][481][0]=96'h7b74;
sos_loop[0].somModel.sram_ptr[7][481]=3;
sos_loop[0].somModel.sram_dat[7][482][0]=96'h117f;
sos_loop[0].somModel.sram_ptr[7][482]=3;
sos_loop[0].somModel.sram_dat[7][483][0]=96'ha024;
sos_loop[0].somModel.sram_ptr[7][483]=3;
sos_loop[0].somModel.sram_dat[7][484][0]=96'hb6cc;
sos_loop[0].somModel.sram_ptr[7][484]=3;
sos_loop[0].somModel.sram_dat[7][485][0]=96'h5a3f;
sos_loop[0].somModel.sram_ptr[7][485]=3;
sos_loop[0].somModel.sram_dat[7][486][0]=96'hbf61;
sos_loop[0].somModel.sram_ptr[7][486]=3;
sos_loop[0].somModel.sram_dat[7][487][0]=96'hc96b;
sos_loop[0].somModel.sram_ptr[7][487]=3;
sos_loop[0].somModel.sram_dat[7][488][0]=96'hc476;
sos_loop[0].somModel.sram_ptr[7][488]=3;
sos_loop[0].somModel.sram_dat[7][489][0]=96'hc029;
sos_loop[0].somModel.sram_ptr[7][489]=3;
sos_loop[0].somModel.sram_dat[7][490][0]=96'h446f;
sos_loop[0].somModel.sram_ptr[7][490]=3;
sos_loop[0].somModel.sram_dat[7][491][0]=96'hc986;
sos_loop[0].somModel.sram_ptr[7][491]=3;
sos_loop[0].somModel.sram_dat[7][492][0]=96'h8bf2;
sos_loop[0].somModel.sram_ptr[7][492]=3;
sos_loop[0].somModel.sram_dat[7][493][0]=96'h190b;
sos_loop[0].somModel.sram_ptr[7][493]=3;
sos_loop[0].somModel.sram_dat[7][494][0]=96'h2afd;
sos_loop[0].somModel.sram_ptr[7][494]=3;
sos_loop[0].somModel.sram_dat[7][495][0]=96'h9aad;
sos_loop[0].somModel.sram_ptr[7][495]=3;
sos_loop[0].somModel.sram_dat[7][496][0]=96'he797;
sos_loop[0].somModel.sram_ptr[7][496]=3;
sos_loop[0].somModel.sram_dat[7][497][0]=96'hc09a;
sos_loop[0].somModel.sram_ptr[7][497]=3;
sos_loop[0].somModel.sram_dat[7][498][0]=96'h671f;
sos_loop[0].somModel.sram_ptr[7][498]=3;
sos_loop[0].somModel.sram_dat[7][499][0]=96'h4c2c;
sos_loop[0].somModel.sram_ptr[7][499]=3;
sos_loop[0].somModel.sram_dat[7][500][0]=96'h3ef1;
sos_loop[0].somModel.sram_ptr[7][500]=3;
sos_loop[0].somModel.sram_dat[7][501][0]=96'hc600;
sos_loop[0].somModel.sram_ptr[7][501]=3;
sos_loop[0].somModel.sram_dat[7][502][0]=96'h6ce5;
sos_loop[0].somModel.sram_ptr[7][502]=3;
sos_loop[0].somModel.sram_dat[7][503][0]=96'h1228;
sos_loop[0].somModel.sram_ptr[7][503]=3;
sos_loop[0].somModel.sram_dat[7][504][0]=96'he80e;
sos_loop[0].somModel.sram_ptr[7][504]=3;
sos_loop[0].somModel.sram_dat[7][505][0]=96'h8dd7;
sos_loop[0].somModel.sram_ptr[7][505]=3;
sos_loop[0].somModel.sram_dat[7][506][0]=96'hd9ff;
sos_loop[0].somModel.sram_ptr[7][506]=3;
sos_loop[0].somModel.sram_dat[7][507][0]=96'h9114;
sos_loop[0].somModel.sram_ptr[7][507]=3;
sos_loop[0].somModel.sram_dat[7][508][0]=96'hfffd;
sos_loop[0].somModel.sram_ptr[7][508]=3;
sos_loop[0].somModel.sram_dat[7][509][0]=96'hfec1;
sos_loop[0].somModel.sram_ptr[7][509]=3;
sos_loop[0].somModel.sram_dat[7][510][0]=96'h157a;
sos_loop[0].somModel.sram_ptr[7][510]=3;
sos_loop[0].somModel.sram_dat[7][511][0]=96'h8698;
sos_loop[0].somModel.sram_ptr[7][511]=3;
sos_loop[0].somModel.sram_dat[7][512][0]=96'h64dd;
sos_loop[0].somModel.sram_ptr[7][512]=3;
sos_loop[0].somModel.sram_dat[7][513][0]=96'h6c7b;
sos_loop[0].somModel.sram_ptr[7][513]=3;
sos_loop[0].somModel.sram_dat[7][514][0]=96'hd6f6;
sos_loop[0].somModel.sram_ptr[7][514]=3;
sos_loop[0].somModel.sram_dat[7][515][0]=96'hd74e;
sos_loop[0].somModel.sram_ptr[7][515]=3;
sos_loop[0].somModel.sram_dat[7][516][0]=96'hd5ca;
sos_loop[0].somModel.sram_ptr[7][516]=3;
sos_loop[0].somModel.sram_dat[7][517][0]=96'h7199;
sos_loop[0].somModel.sram_ptr[7][517]=3;
sos_loop[0].somModel.sram_dat[7][518][0]=96'h5167;
sos_loop[0].somModel.sram_ptr[7][518]=3;
sos_loop[0].somModel.sram_dat[7][519][0]=96'h2b74;
sos_loop[0].somModel.sram_ptr[7][519]=3;
sos_loop[0].somModel.sram_dat[7][520][0]=96'h418b;
sos_loop[0].somModel.sram_ptr[7][520]=3;
sos_loop[0].somModel.sram_dat[7][521][0]=96'h4e9a;
sos_loop[0].somModel.sram_ptr[7][521]=3;
sos_loop[0].somModel.sram_dat[7][522][0]=96'h8692;
sos_loop[0].somModel.sram_ptr[7][522]=3;
sos_loop[0].somModel.sram_dat[7][523][0]=96'hc6e0;
sos_loop[0].somModel.sram_ptr[7][523]=3;
sos_loop[0].somModel.sram_dat[7][524][0]=96'h1f44;
sos_loop[0].somModel.sram_ptr[7][524]=3;
sos_loop[0].somModel.sram_dat[7][525][0]=96'h75a0;
sos_loop[0].somModel.sram_ptr[7][525]=3;
sos_loop[0].somModel.sram_dat[7][526][0]=96'h3793;
sos_loop[0].somModel.sram_ptr[7][526]=3;
sos_loop[0].somModel.sram_dat[7][527][0]=96'h6365;
sos_loop[0].somModel.sram_ptr[7][527]=3;
sos_loop[0].somModel.sram_dat[7][528][0]=96'hee99;
sos_loop[0].somModel.sram_ptr[7][528]=3;
sos_loop[0].somModel.sram_dat[7][529][0]=96'hac5;
sos_loop[0].somModel.sram_ptr[7][529]=3;
sos_loop[0].somModel.sram_dat[7][530][0]=96'h6b09;
sos_loop[0].somModel.sram_ptr[7][530]=3;
sos_loop[0].somModel.sram_dat[7][531][0]=96'h54d0;
sos_loop[0].somModel.sram_ptr[7][531]=3;
sos_loop[0].somModel.sram_dat[7][532][0]=96'hb98d;
sos_loop[0].somModel.sram_ptr[7][532]=3;
sos_loop[0].somModel.sram_dat[7][533][0]=96'hd586;
sos_loop[0].somModel.sram_ptr[7][533]=3;
sos_loop[0].somModel.sram_dat[7][534][0]=96'h4cc3;
sos_loop[0].somModel.sram_ptr[7][534]=3;
sos_loop[0].somModel.sram_dat[7][535][0]=96'hc26c;
sos_loop[0].somModel.sram_ptr[7][535]=3;
sos_loop[0].somModel.sram_dat[7][536][0]=96'hf681;
sos_loop[0].somModel.sram_ptr[7][536]=3;
sos_loop[0].somModel.sram_dat[7][537][0]=96'hf0c9;
sos_loop[0].somModel.sram_ptr[7][537]=3;
sos_loop[0].somModel.sram_dat[7][538][0]=96'hbe02;
sos_loop[0].somModel.sram_ptr[7][538]=3;
sos_loop[0].somModel.sram_dat[7][539][0]=96'h5eb8;
sos_loop[0].somModel.sram_ptr[7][539]=3;
sos_loop[0].somModel.sram_dat[7][540][0]=96'h4c1e;
sos_loop[0].somModel.sram_ptr[7][540]=3;
sos_loop[0].somModel.sram_dat[7][541][0]=96'hc52a;
sos_loop[0].somModel.sram_ptr[7][541]=3;
sos_loop[0].somModel.sram_dat[7][542][0]=96'h93c;
sos_loop[0].somModel.sram_ptr[7][542]=3;
sos_loop[0].somModel.sram_dat[7][543][0]=96'hd07f;
sos_loop[0].somModel.sram_ptr[7][543]=3;
sos_loop[0].somModel.sram_dat[7][544][0]=96'hd767;
sos_loop[0].somModel.sram_ptr[7][544]=3;
sos_loop[0].somModel.sram_dat[7][545][0]=96'h29db;
sos_loop[0].somModel.sram_ptr[7][545]=3;
sos_loop[0].somModel.sram_dat[7][546][0]=96'h2546;
sos_loop[0].somModel.sram_ptr[7][546]=3;
sos_loop[0].somModel.sram_dat[7][547][0]=96'h12d9;
sos_loop[0].somModel.sram_ptr[7][547]=3;
sos_loop[0].somModel.sram_dat[7][548][0]=96'hff67;
sos_loop[0].somModel.sram_ptr[7][548]=3;
sos_loop[0].somModel.sram_dat[7][549][0]=96'hda73;
sos_loop[0].somModel.sram_ptr[7][549]=3;
sos_loop[0].somModel.sram_dat[7][550][0]=96'hb6d;
sos_loop[0].somModel.sram_ptr[7][550]=3;
sos_loop[0].somModel.sram_dat[7][551][0]=96'hf5b5;
sos_loop[0].somModel.sram_ptr[7][551]=3;
sos_loop[0].somModel.sram_dat[7][552][0]=96'h6e7;
sos_loop[0].somModel.sram_ptr[7][552]=3;
sos_loop[0].somModel.sram_dat[7][553][0]=96'hd236;
sos_loop[0].somModel.sram_ptr[7][553]=3;
sos_loop[0].somModel.sram_dat[7][554][0]=96'hb505;
sos_loop[0].somModel.sram_ptr[7][554]=3;
sos_loop[0].somModel.sram_dat[7][555][0]=96'h7813;
sos_loop[0].somModel.sram_ptr[7][555]=3;
sos_loop[0].somModel.sram_dat[7][556][0]=96'h199a;
sos_loop[0].somModel.sram_ptr[7][556]=3;
sos_loop[0].somModel.sram_dat[7][557][0]=96'h1e9d;
sos_loop[0].somModel.sram_ptr[7][557]=3;
sos_loop[0].somModel.sram_dat[7][558][0]=96'h8438;
sos_loop[0].somModel.sram_ptr[7][558]=3;
sos_loop[0].somModel.sram_dat[7][559][0]=96'h853c;
sos_loop[0].somModel.sram_ptr[7][559]=3;
sos_loop[0].somModel.sram_dat[7][560][0]=96'hfa90;
sos_loop[0].somModel.sram_ptr[7][560]=3;
sos_loop[0].somModel.sram_dat[7][561][0]=96'h91d3;
sos_loop[0].somModel.sram_ptr[7][561]=3;
sos_loop[0].somModel.sram_dat[7][562][0]=96'h9871;
sos_loop[0].somModel.sram_ptr[7][562]=3;
sos_loop[0].somModel.sram_dat[7][563][0]=96'hf155;
sos_loop[0].somModel.sram_ptr[7][563]=3;
sos_loop[0].somModel.sram_dat[7][564][0]=96'hec3;
sos_loop[0].somModel.sram_ptr[7][564]=3;
sos_loop[0].somModel.sram_dat[7][565][0]=96'h240;
sos_loop[0].somModel.sram_ptr[7][565]=3;
sos_loop[0].somModel.sram_dat[7][566][0]=96'hc7bf;
sos_loop[0].somModel.sram_ptr[7][566]=3;
sos_loop[0].somModel.sram_dat[7][567][0]=96'h3579;
sos_loop[0].somModel.sram_ptr[7][567]=3;
sos_loop[0].somModel.sram_dat[7][568][0]=96'h6f16;
sos_loop[0].somModel.sram_ptr[7][568]=3;
sos_loop[0].somModel.sram_dat[7][569][0]=96'h2fbd;
sos_loop[0].somModel.sram_ptr[7][569]=3;
sos_loop[0].somModel.sram_dat[7][570][0]=96'h376f;
sos_loop[0].somModel.sram_ptr[7][570]=3;
sos_loop[0].somModel.sram_dat[7][571][0]=96'h8129;
sos_loop[0].somModel.sram_ptr[7][571]=3;
sos_loop[0].somModel.sram_dat[7][572][0]=96'hcb9c;
sos_loop[0].somModel.sram_ptr[7][572]=3;
sos_loop[0].somModel.sram_dat[7][573][0]=96'h8b5a;
sos_loop[0].somModel.sram_ptr[7][573]=3;
sos_loop[0].somModel.sram_dat[7][574][0]=96'hc137;
sos_loop[0].somModel.sram_ptr[7][574]=3;
sos_loop[0].somModel.sram_dat[7][575][0]=96'h16b5;
sos_loop[0].somModel.sram_ptr[7][575]=3;
sos_loop[0].somModel.sram_dat[7][576][0]=96'h9006;
sos_loop[0].somModel.sram_ptr[7][576]=3;
sos_loop[0].somModel.sram_dat[7][577][0]=96'h24fd;
sos_loop[0].somModel.sram_ptr[7][577]=3;
sos_loop[0].somModel.sram_dat[7][578][0]=96'h38c7;
sos_loop[0].somModel.sram_ptr[7][578]=3;
sos_loop[0].somModel.sram_dat[7][579][0]=96'hf065;
sos_loop[0].somModel.sram_ptr[7][579]=3;
sos_loop[0].somModel.sram_dat[7][580][0]=96'hd149;
sos_loop[0].somModel.sram_ptr[7][580]=3;
sos_loop[0].somModel.sram_dat[7][581][0]=96'hf573;
sos_loop[0].somModel.sram_ptr[7][581]=3;
sos_loop[0].somModel.sram_dat[7][582][0]=96'ha7e5;
sos_loop[0].somModel.sram_ptr[7][582]=3;
sos_loop[0].somModel.sram_dat[7][583][0]=96'hc110;
sos_loop[0].somModel.sram_ptr[7][583]=3;
sos_loop[0].somModel.sram_dat[7][584][0]=96'h6859;
sos_loop[0].somModel.sram_ptr[7][584]=3;
sos_loop[0].somModel.sram_dat[7][585][0]=96'h66bb;
sos_loop[0].somModel.sram_ptr[7][585]=3;
sos_loop[0].somModel.sram_dat[7][586][0]=96'h6dc2;
sos_loop[0].somModel.sram_ptr[7][586]=3;
sos_loop[0].somModel.sram_dat[7][587][0]=96'hfce5;
sos_loop[0].somModel.sram_ptr[7][587]=3;
sos_loop[0].somModel.sram_dat[7][588][0]=96'h89f3;
sos_loop[0].somModel.sram_ptr[7][588]=3;
sos_loop[0].somModel.sram_dat[7][589][0]=96'h188f;
sos_loop[0].somModel.sram_ptr[7][589]=3;
sos_loop[0].somModel.sram_dat[7][590][0]=96'hc76;
sos_loop[0].somModel.sram_ptr[7][590]=3;
sos_loop[0].somModel.sram_dat[7][591][0]=96'hd66;
sos_loop[0].somModel.sram_ptr[7][591]=3;
sos_loop[0].somModel.sram_dat[7][592][0]=96'h8a86;
sos_loop[0].somModel.sram_ptr[7][592]=3;
sos_loop[0].somModel.sram_dat[7][593][0]=96'h2056;
sos_loop[0].somModel.sram_ptr[7][593]=3;
sos_loop[0].somModel.sram_dat[7][594][0]=96'hc598;
sos_loop[0].somModel.sram_ptr[7][594]=3;
sos_loop[0].somModel.sram_dat[7][595][0]=96'h1cb6;
sos_loop[0].somModel.sram_ptr[7][595]=3;
sos_loop[0].somModel.sram_dat[7][596][0]=96'h79c6;
sos_loop[0].somModel.sram_ptr[7][596]=3;
sos_loop[0].somModel.sram_dat[7][597][0]=96'h7621;
sos_loop[0].somModel.sram_ptr[7][597]=3;
sos_loop[0].somModel.sram_dat[7][598][0]=96'hbd5d;
sos_loop[0].somModel.sram_ptr[7][598]=3;
sos_loop[0].somModel.sram_dat[7][599][0]=96'h80e8;
sos_loop[0].somModel.sram_ptr[7][599]=3;
sos_loop[0].somModel.sram_dat[7][600][0]=96'h581f;
sos_loop[0].somModel.sram_ptr[7][600]=3;
sos_loop[0].somModel.sram_dat[7][601][0]=96'hc915;
sos_loop[0].somModel.sram_ptr[7][601]=3;
sos_loop[0].somModel.sram_dat[7][602][0]=96'h1142;
sos_loop[0].somModel.sram_ptr[7][602]=3;
sos_loop[0].somModel.sram_dat[7][603][0]=96'h39df;
sos_loop[0].somModel.sram_ptr[7][603]=3;
sos_loop[0].somModel.sram_dat[7][604][0]=96'h55cc;
sos_loop[0].somModel.sram_ptr[7][604]=3;
sos_loop[0].somModel.sram_dat[7][605][0]=96'hf2a1;
sos_loop[0].somModel.sram_ptr[7][605]=3;
sos_loop[0].somModel.sram_dat[7][606][0]=96'hfa13;
sos_loop[0].somModel.sram_ptr[7][606]=3;
sos_loop[0].somModel.sram_dat[7][607][0]=96'h4c4;
sos_loop[0].somModel.sram_ptr[7][607]=3;
sos_loop[0].somModel.sram_dat[7][608][0]=96'haa67;
sos_loop[0].somModel.sram_ptr[7][608]=3;
sos_loop[0].somModel.sram_dat[7][609][0]=96'h187a;
sos_loop[0].somModel.sram_ptr[7][609]=3;
sos_loop[0].somModel.sram_dat[7][610][0]=96'h8437;
sos_loop[0].somModel.sram_ptr[7][610]=3;
sos_loop[0].somModel.sram_dat[7][611][0]=96'hfaf;
sos_loop[0].somModel.sram_ptr[7][611]=3;
sos_loop[0].somModel.sram_dat[7][612][0]=96'h10bb;
sos_loop[0].somModel.sram_ptr[7][612]=3;
sos_loop[0].somModel.sram_dat[7][613][0]=96'hc03c;
sos_loop[0].somModel.sram_ptr[7][613]=3;
sos_loop[0].somModel.sram_dat[7][614][0]=96'ha17d;
sos_loop[0].somModel.sram_ptr[7][614]=3;
sos_loop[0].somModel.sram_dat[7][615][0]=96'ha172;
sos_loop[0].somModel.sram_ptr[7][615]=3;
sos_loop[0].somModel.sram_dat[7][616][0]=96'h36c5;
sos_loop[0].somModel.sram_ptr[7][616]=3;
sos_loop[0].somModel.sram_dat[7][617][0]=96'h344d;
sos_loop[0].somModel.sram_ptr[7][617]=3;
sos_loop[0].somModel.sram_dat[7][618][0]=96'h4e82;
sos_loop[0].somModel.sram_ptr[7][618]=3;
sos_loop[0].somModel.sram_dat[7][619][0]=96'he473;
sos_loop[0].somModel.sram_ptr[7][619]=3;
sos_loop[0].somModel.sram_dat[7][620][0]=96'h4bfd;
sos_loop[0].somModel.sram_ptr[7][620]=3;
sos_loop[0].somModel.sram_dat[7][621][0]=96'hd436;
sos_loop[0].somModel.sram_ptr[7][621]=3;
sos_loop[0].somModel.sram_dat[7][622][0]=96'h33a7;
sos_loop[0].somModel.sram_ptr[7][622]=3;
sos_loop[0].somModel.sram_dat[7][623][0]=96'he4bf;
sos_loop[0].somModel.sram_ptr[7][623]=3;
sos_loop[0].somModel.sram_dat[7][624][0]=96'h4c20;
sos_loop[0].somModel.sram_ptr[7][624]=3;
sos_loop[0].somModel.sram_dat[7][625][0]=96'hc7cc;
sos_loop[0].somModel.sram_ptr[7][625]=3;
sos_loop[0].somModel.sram_dat[7][626][0]=96'h2ff0;
sos_loop[0].somModel.sram_ptr[7][626]=3;
sos_loop[0].somModel.sram_dat[7][627][0]=96'h33c8;
sos_loop[0].somModel.sram_ptr[7][627]=3;
sos_loop[0].somModel.sram_dat[7][628][0]=96'h40c4;
sos_loop[0].somModel.sram_ptr[7][628]=3;
sos_loop[0].somModel.sram_dat[7][629][0]=96'h64a9;
sos_loop[0].somModel.sram_ptr[7][629]=3;
sos_loop[0].somModel.sram_dat[7][630][0]=96'h78d;
sos_loop[0].somModel.sram_ptr[7][630]=3;
sos_loop[0].somModel.sram_dat[7][631][0]=96'ha2d3;
sos_loop[0].somModel.sram_ptr[7][631]=3;
sos_loop[0].somModel.sram_dat[7][632][0]=96'h3326;
sos_loop[0].somModel.sram_ptr[7][632]=3;
sos_loop[0].somModel.sram_dat[7][633][0]=96'hdbf9;
sos_loop[0].somModel.sram_ptr[7][633]=3;
sos_loop[0].somModel.sram_dat[7][634][0]=96'h907a;
sos_loop[0].somModel.sram_ptr[7][634]=3;
sos_loop[0].somModel.sram_dat[7][635][0]=96'he187;
sos_loop[0].somModel.sram_ptr[7][635]=3;
sos_loop[0].somModel.sram_dat[7][636][0]=96'h1c66;
sos_loop[0].somModel.sram_ptr[7][636]=3;
sos_loop[0].somModel.sram_dat[7][637][0]=96'hf67e;
sos_loop[0].somModel.sram_ptr[7][637]=3;
sos_loop[0].somModel.sram_dat[7][638][0]=96'h4aa1;
sos_loop[0].somModel.sram_ptr[7][638]=3;
sos_loop[0].somModel.sram_dat[7][639][0]=96'hfd6b;
sos_loop[0].somModel.sram_ptr[7][639]=3;
sos_loop[0].somModel.sram_dat[7][640][0]=96'hb65b;
sos_loop[0].somModel.sram_ptr[7][640]=3;
sos_loop[0].somModel.sram_dat[7][641][0]=96'h50f8;
sos_loop[0].somModel.sram_ptr[7][641]=3;
sos_loop[0].somModel.sram_dat[7][642][0]=96'hee03;
sos_loop[0].somModel.sram_ptr[7][642]=3;
sos_loop[0].somModel.sram_dat[7][643][0]=96'hbf2d;
sos_loop[0].somModel.sram_ptr[7][643]=3;
sos_loop[0].somModel.sram_dat[7][644][0]=96'h5809;
sos_loop[0].somModel.sram_ptr[7][644]=3;
sos_loop[0].somModel.sram_dat[7][645][0]=96'he9a7;
sos_loop[0].somModel.sram_ptr[7][645]=3;
sos_loop[0].somModel.sram_dat[7][646][0]=96'hf3f3;
sos_loop[0].somModel.sram_ptr[7][646]=3;
sos_loop[0].somModel.sram_dat[7][647][0]=96'h8ce2;
sos_loop[0].somModel.sram_ptr[7][647]=3;
sos_loop[0].somModel.sram_dat[7][648][0]=96'hc953;
sos_loop[0].somModel.sram_ptr[7][648]=3;
sos_loop[0].somModel.sram_dat[7][649][0]=96'hb0d;
sos_loop[0].somModel.sram_ptr[7][649]=3;
sos_loop[0].somModel.sram_dat[7][650][0]=96'h623b;
sos_loop[0].somModel.sram_ptr[7][650]=3;
sos_loop[0].somModel.sram_dat[7][651][0]=96'ha57a;
sos_loop[0].somModel.sram_ptr[7][651]=3;
sos_loop[0].somModel.sram_dat[7][652][0]=96'hbbfd;
sos_loop[0].somModel.sram_ptr[7][652]=3;
sos_loop[0].somModel.sram_dat[7][653][0]=96'hcd5;
sos_loop[0].somModel.sram_ptr[7][653]=3;
sos_loop[0].somModel.sram_dat[7][654][0]=96'h7d9;
sos_loop[0].somModel.sram_ptr[7][654]=3;
sos_loop[0].somModel.sram_dat[7][655][0]=96'hd5b7;
sos_loop[0].somModel.sram_ptr[7][655]=3;
sos_loop[0].somModel.sram_dat[7][656][0]=96'hc765;
sos_loop[0].somModel.sram_ptr[7][656]=3;
sos_loop[0].somModel.sram_dat[7][657][0]=96'haf71;
sos_loop[0].somModel.sram_ptr[7][657]=3;
sos_loop[0].somModel.sram_dat[7][658][0]=96'he0e2;
sos_loop[0].somModel.sram_ptr[7][658]=3;
sos_loop[0].somModel.sram_dat[7][659][0]=96'heab4;
sos_loop[0].somModel.sram_ptr[7][659]=3;
sos_loop[0].somModel.sram_dat[7][660][0]=96'hb006;
sos_loop[0].somModel.sram_ptr[7][660]=3;
sos_loop[0].somModel.sram_dat[7][661][0]=96'ha268;
sos_loop[0].somModel.sram_ptr[7][661]=3;
sos_loop[0].somModel.sram_dat[7][662][0]=96'h2e18;
sos_loop[0].somModel.sram_ptr[7][662]=3;
sos_loop[0].somModel.sram_dat[7][663][0]=96'h8f7d;
sos_loop[0].somModel.sram_ptr[7][663]=3;
sos_loop[0].somModel.sram_dat[7][664][0]=96'hb733;
sos_loop[0].somModel.sram_ptr[7][664]=3;
sos_loop[0].somModel.sram_dat[7][665][0]=96'h7454;
sos_loop[0].somModel.sram_ptr[7][665]=3;
sos_loop[0].somModel.sram_dat[7][666][0]=96'h651;
sos_loop[0].somModel.sram_ptr[7][666]=3;
sos_loop[0].somModel.sram_dat[7][667][0]=96'h21c7;
sos_loop[0].somModel.sram_ptr[7][667]=3;
sos_loop[0].somModel.sram_dat[7][668][0]=96'hf615;
sos_loop[0].somModel.sram_ptr[7][668]=3;
sos_loop[0].somModel.sram_dat[7][669][0]=96'hd932;
sos_loop[0].somModel.sram_ptr[7][669]=3;
sos_loop[0].somModel.sram_dat[7][670][0]=96'hdc24;
sos_loop[0].somModel.sram_ptr[7][670]=3;
sos_loop[0].somModel.sram_dat[7][671][0]=96'h6b3b;
sos_loop[0].somModel.sram_ptr[7][671]=3;
sos_loop[0].somModel.sram_dat[7][672][0]=96'ha575;
sos_loop[0].somModel.sram_ptr[7][672]=3;
sos_loop[0].somModel.sram_dat[7][673][0]=96'h7f07;
sos_loop[0].somModel.sram_ptr[7][673]=3;
sos_loop[0].somModel.sram_dat[7][674][0]=96'hbb77;
sos_loop[0].somModel.sram_ptr[7][674]=3;
sos_loop[0].somModel.sram_dat[7][675][0]=96'h4308;
sos_loop[0].somModel.sram_ptr[7][675]=3;
sos_loop[0].somModel.sram_dat[7][676][0]=96'h901d;
sos_loop[0].somModel.sram_ptr[7][676]=3;
sos_loop[0].somModel.sram_dat[7][677][0]=96'h2f04;
sos_loop[0].somModel.sram_ptr[7][677]=3;
sos_loop[0].somModel.sram_dat[7][678][0]=96'h672;
sos_loop[0].somModel.sram_ptr[7][678]=3;
sos_loop[0].somModel.sram_dat[7][679][0]=96'h4440;
sos_loop[0].somModel.sram_ptr[7][679]=3;
sos_loop[0].somModel.sram_dat[7][680][0]=96'h222;
sos_loop[0].somModel.sram_ptr[7][680]=3;
sos_loop[0].somModel.sram_dat[7][681][0]=96'h208f;
sos_loop[0].somModel.sram_ptr[7][681]=3;
sos_loop[0].somModel.sram_dat[7][682][0]=96'hb0a7;
sos_loop[0].somModel.sram_ptr[7][682]=3;
sos_loop[0].somModel.sram_dat[7][683][0]=96'h1a32;
sos_loop[0].somModel.sram_ptr[7][683]=3;
sos_loop[0].somModel.sram_dat[7][684][0]=96'hb3cd;
sos_loop[0].somModel.sram_ptr[7][684]=3;
sos_loop[0].somModel.sram_dat[7][685][0]=96'hcef3;
sos_loop[0].somModel.sram_ptr[7][685]=3;
sos_loop[0].somModel.sram_dat[7][686][0]=96'h5f33;
sos_loop[0].somModel.sram_ptr[7][686]=3;
sos_loop[0].somModel.sram_dat[7][687][0]=96'h5003;
sos_loop[0].somModel.sram_ptr[7][687]=3;
sos_loop[0].somModel.sram_dat[7][688][0]=96'h2cb3;
sos_loop[0].somModel.sram_ptr[7][688]=3;
sos_loop[0].somModel.sram_dat[7][689][0]=96'hf670;
sos_loop[0].somModel.sram_ptr[7][689]=3;
sos_loop[0].somModel.sram_dat[7][690][0]=96'hb8be;
sos_loop[0].somModel.sram_ptr[7][690]=3;
sos_loop[0].somModel.sram_dat[7][691][0]=96'h254b;
sos_loop[0].somModel.sram_ptr[7][691]=3;
sos_loop[0].somModel.sram_dat[7][692][0]=96'hb525;
sos_loop[0].somModel.sram_ptr[7][692]=3;
sos_loop[0].somModel.sram_dat[7][693][0]=96'h9a07;
sos_loop[0].somModel.sram_ptr[7][693]=3;
sos_loop[0].somModel.sram_dat[7][694][0]=96'haf14;
sos_loop[0].somModel.sram_ptr[7][694]=3;
sos_loop[0].somModel.sram_dat[7][695][0]=96'h759e;
sos_loop[0].somModel.sram_ptr[7][695]=3;
sos_loop[0].somModel.sram_dat[7][696][0]=96'hd9b5;
sos_loop[0].somModel.sram_ptr[7][696]=3;
sos_loop[0].somModel.sram_dat[7][697][0]=96'h2612;
sos_loop[0].somModel.sram_ptr[7][697]=3;
sos_loop[0].somModel.sram_dat[7][698][0]=96'he49c;
sos_loop[0].somModel.sram_ptr[7][698]=3;
sos_loop[0].somModel.sram_dat[7][699][0]=96'hfc4a;
sos_loop[0].somModel.sram_ptr[7][699]=3;
sos_loop[0].somModel.sram_dat[7][700][0]=96'hd6fd;
sos_loop[0].somModel.sram_ptr[7][700]=3;
sos_loop[0].somModel.cfg_tbl_sel[7] = 7;
sos_loop[0].somModel.cfg_dat_sel[7] = 2;
sos_loop[0].somModel.cfg_dat_vld[7] = 1;
sos_loop[0].somModel.cfg_miss_ptr[7] = 0;
end