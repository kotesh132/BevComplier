add_config_entry(0, 32'hc0, 2, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000083);
add_config_entry(0, 32'hc2, 2, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000045);
add_config_entry(0, 32'hc4, 2, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080000087);
add_config_entry(0, 32'hc6, 2, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000209);
add_config_entry(0, 32'hc8, 2, 512'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040000040b);
add_config_entry(0, 32'hca, 2, 512'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000004d);
add_config_entry(0, 32'hcc, 2, 512'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010f);
add_config_entry(0, 32'h80, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
add_config_entry(0, 32'h81, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008);
add_config_entry(0, 32'h82, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010);
add_config_entry(0, 32'h83, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018);
add_config_entry(0, 32'h84, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020);
add_config_entry(0, 32'h85, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000028);
add_config_entry(0, 32'h86, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000030);
add_config_entry(0, 32'h87, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
add_config_entry(0, 32'h88, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
add_config_entry(0, 32'h89, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
add_config_entry(0, 32'h8a, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
add_config_entry(0, 32'h8b, 1, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
add_config_entry(0, 32'ha0, 2, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009);
add_config_entry(0, 32'ha2, 2, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000005);
add_config_entry(0, 32'ha4, 2, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000081);
add_config_entry(0, 32'ha6, 2, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000011);
add_config_entry(0, 32'ha8, 2, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000400000101);
add_config_entry(0, 32'haa, 2, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000600000021);
add_config_entry(0, 32'hac, 2, 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000800000041);
add_config_entry(0, 32'h40, 3, 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007fe000200000000021);
add_config_entry(0, 32'h43, 3, 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007fe000200800000011);
add_config_entry(0, 32'h46, 3, 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007fe000200000000201);
add_config_entry(0, 32'h49, 3, 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007fe000200800000041);
add_config_entry(0, 32'h4c, 3, 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007fe000201000000401);
add_config_entry(0, 32'h4f, 3, 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007fe000201800000081);
add_config_entry(0, 32'h52, 3, 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007fe000202000000101);
