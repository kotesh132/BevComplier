initial begin
@(posedge clk);
@(negedge rst);
@(posedge clk);
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[1] = 80'h9b2571c7073c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[1] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[2] = 80'hede35ed4bae4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[2] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[3] = 80'hd835b1486b13;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[3] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[4] = 80'hbe3dd6d14071;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[4] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[5] = 80'h88e0f6aa248a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[5] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[6] = 80'hf3012b605570;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[6] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[7] = 80'he16202381133;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[7] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[8] = 80'hf16aa927fb4a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[8] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[9] = 80'h458011f44fab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[9] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[10] = 80'h6b5603b74017;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[10] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[11] = 80'h9867863b5169;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[11] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[12] = 80'h7d563611e661;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[12] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[13] = 80'h9a388934f048;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[13] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[14] = 80'he7d208135786;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[14] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[15] = 80'h1d236be012e4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[15] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[16] = 80'h4816ad6457a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[16] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[17] = 80'hb7fcfacfa875;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[17] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[18] = 80'hacdaf0aca7c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[18] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[19] = 80'h272061475aea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[19] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[20] = 80'hed5c1ad98d27;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[20] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[21] = 80'h5137add3842;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[21] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[22] = 80'h77c13eb8f0bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[22] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[23] = 80'h64dec849f297;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[23] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[24] = 80'h52815aaa0e76;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[24] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[25] = 80'h36c627639625;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[25] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[26] = 80'hadfa0e35ab63;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[26] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[27] = 80'hde873f211f1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[27] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[28] = 80'h7c056a29eb06;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[28] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[29] = 80'hb17370ad5889;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[29] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[30] = 80'h3c16a3b80a77;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[30] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[31] = 80'hfdc75e2fe46f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[31] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[32] = 80'hb514aca9a7ea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[32] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[33] = 80'hff4fc0b5dd4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[33] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[34] = 80'h4fa3edb32414;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[34] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[35] = 80'ha7a0a91df8ba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[35] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[36] = 80'hf1dccb540bd9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[36] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[37] = 80'hdb32f0046c0d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[37] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[38] = 80'h5be7f8e59bc2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[38] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[39] = 80'h56ae936d2b74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[39] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[40] = 80'h21237dd3755f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[40] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[41] = 80'ha6839f79036b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[41] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[42] = 80'h5e54e001a27;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[42] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[43] = 80'h2dfc19bbb79a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[43] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[44] = 80'h7da11a068ee0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[44] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[45] = 80'h7b392b497f6e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[45] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[46] = 80'h6c0398426174;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[46] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[47] = 80'h7b724903d7a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[47] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[48] = 80'h7e2e109e6271;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[48] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[49] = 80'h70b0857e229f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[49] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[50] = 80'h276af0ce7d95;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[50] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[51] = 80'h977c2662d661;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[51] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[52] = 80'h6c110a6ebb5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[52] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[53] = 80'h7100f4f63c98;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[53] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[54] = 80'hdee6b07e350;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[54] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[55] = 80'h73f1bab9b30b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[55] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[56] = 80'h45a7a7cd7c56;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[56] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[57] = 80'h5c2982129594;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[57] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[58] = 80'h24f31697e85b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[58] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[59] = 80'h1217e5938719;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[59] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[60] = 80'hd7165d2854bd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[60] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[61] = 80'ha943cd77303b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[61] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[62] = 80'heb90c7477f53;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[62] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[63] = 80'h445c3e0895fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[63] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[64] = 80'hb312060a0eef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[64] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[65] = 80'hcc66a816d743;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[65] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[66] = 80'hb3497a7141e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[66] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[67] = 80'h822765751942;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[67] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[68] = 80'h199ff6767d07;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[68] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[69] = 80'hd15a97c2415f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[69] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[70] = 80'he029b33bdf0c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[70] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[71] = 80'h516f120d3a96;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[71] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[72] = 80'h4e9aec95e85c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[72] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[73] = 80'hd172c141c22a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[73] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[74] = 80'h73147f2a5ee0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[74] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[75] = 80'hfbb8275391e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[75] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[76] = 80'h65fdd1b8aab4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[76] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[77] = 80'hf1874d4b4c76;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[77] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[78] = 80'h6cd16dcc4a33;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[78] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[79] = 80'hd96441dc2078;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[79] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[80] = 80'hc319811fd277;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[80] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[81] = 80'h8a0471dd6d11;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[81] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[82] = 80'hf394863f8076;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[82] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[83] = 80'h5b121b7039e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[83] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[84] = 80'heafeaba615dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[84] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[85] = 80'hc10aef68e81f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[85] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[86] = 80'hb4285b984022;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[86] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[87] = 80'h8264ffadb985;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[87] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[88] = 80'ha5638ebc9ea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[88] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[89] = 80'hc025ca05681b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[89] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[90] = 80'h69fc597ace55;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[90] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[91] = 80'h92d13ceb35ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[91] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[92] = 80'hd92c798e2da4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[92] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[93] = 80'hef44bbde26b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[93] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[94] = 80'h4a7bde16a1b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[94] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[95] = 80'h9cef75742606;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[95] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[96] = 80'hbc689291a89e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[96] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[97] = 80'hecad85584eac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[97] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[98] = 80'h2596ab0bd4ef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[98] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[99] = 80'hafb0bcd5f28c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[99] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[100] = 80'h588ea274f953;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[100] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[101] = 80'ha7391453de54;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[101] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[102] = 80'hfdbcbd10e033;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[102] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[103] = 80'h719cfa2767c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[103] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[104] = 80'ha3ef35e42c33;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[104] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[105] = 80'hc4c69a60a71a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[105] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[106] = 80'h3a3a7b0a793b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[106] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[107] = 80'hcfa4b3cac05c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[107] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[108] = 80'h5599e50df8a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[108] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[109] = 80'h3a0f6debddd0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[109] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[110] = 80'h9f11ab78573a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[110] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[111] = 80'hd608068e6320;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[111] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[112] = 80'hd862045cf75f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[112] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[113] = 80'h6cae027bae23;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[113] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[114] = 80'he2a567e44491;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[114] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[115] = 80'h72c9f8b64ee2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[115] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[116] = 80'h408440fab4cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[116] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[117] = 80'h4309898b60f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[117] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[118] = 80'h115a7eb75e3a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[118] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[119] = 80'h37178729e67f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[119] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[120] = 80'hfb424524db25;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[120] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[121] = 80'h361984d7eb12;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[121] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[122] = 80'h927e86180bf1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[122] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[123] = 80'h6a2879654a57;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[123] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[124] = 80'h641b343f80f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[124] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[125] = 80'h93991f1d7362;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[125] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[126] = 80'h15e87559900d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[126] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[127] = 80'h5d613c992175;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[127] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[128] = 80'h899161eca21b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[128] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[129] = 80'h4a353e6fdb65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[129] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[130] = 80'h6d2289d6b1b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[130] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[131] = 80'h63d6892f4cbd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[131] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[132] = 80'hec516e56e38;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[132] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[133] = 80'hf6d75e867538;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[133] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[134] = 80'hf8103fe52fca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[134] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[135] = 80'h3721758992ed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[135] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[136] = 80'hc7a4b46ded9a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[136] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[137] = 80'h8261693eedaf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[137] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[138] = 80'h3a70bd4ccb71;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[138] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[139] = 80'hdc3e4883a653;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[139] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[140] = 80'h6bb7508ac2dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[140] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[141] = 80'h873638a207ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[141] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[142] = 80'h4732c91bc5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[142] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[143] = 80'h3fd9b4c00a99;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[143] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[144] = 80'h859aa75fc399;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[144] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[145] = 80'h78ba5e9eee08;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[145] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[146] = 80'hdbd3b819af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[146] = 80'hffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[147] = 80'h80957200a77;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[147] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[148] = 80'had807c006574;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[148] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[149] = 80'hb25671eb1928;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[149] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[150] = 80'hcd733d038007;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[150] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[151] = 80'h5a808481d4f8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[151] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[152] = 80'he5270474bc3d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[152] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[153] = 80'h43c133e30238;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[153] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[154] = 80'hda06327c0fb6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[154] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[155] = 80'hf44aa55e8d5b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[155] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[156] = 80'hd108767b16e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[156] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[157] = 80'h45b722c61027;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[157] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[158] = 80'ha633db8c75b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[158] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[159] = 80'hf2d4b44fd6dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[159] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[160] = 80'haffaa97c08bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[160] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[161] = 80'h3db1f6e4e6a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[161] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[162] = 80'hcc8499d91df3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[162] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[163] = 80'hbde381c08689;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[163] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[164] = 80'h4903fd0700cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[164] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[165] = 80'h1af8bbb7c7be;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[165] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[166] = 80'hd7cd2a4ee374;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[166] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[167] = 80'h648e675ea632;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[167] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[168] = 80'h2ab6d3cad9b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[168] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[169] = 80'h5f26b6f13520;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[169] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[170] = 80'ha96772107053;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[170] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[171] = 80'hfd5134dc543a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[171] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[172] = 80'hf9e15e388cda;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[172] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[173] = 80'h37ad0dd04d1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[173] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[174] = 80'h24ed9e62765c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[174] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[175] = 80'hdeaa2a8e2c76;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[175] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[176] = 80'h9afd8ccdf0d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[176] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[177] = 80'hdfba92cc34c0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[177] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[178] = 80'h1d1b77568814;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[178] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[179] = 80'hc138abed4b17;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[179] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[180] = 80'h38fe88806ab3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[180] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[181] = 80'hf4a91c35928f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[181] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[182] = 80'h53d53e8897d5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[182] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[183] = 80'h91213c03913d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[183] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[184] = 80'h39beec93c1a6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[184] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[185] = 80'hb842fcc92642;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[185] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[186] = 80'h5350a885c6e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[186] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[187] = 80'h3a60895d3611;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[187] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[188] = 80'h3958522de12b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[188] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[189] = 80'h8379dd2f10a6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[189] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[190] = 80'h719a6a66e65a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[190] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[191] = 80'h151b0bccc299;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[191] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[192] = 80'h60a3a0ebb851;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[192] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[193] = 80'hceeb751d2978;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[193] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[194] = 80'h6799c24bb3b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[194] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[195] = 80'h56badc0db157;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[195] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[196] = 80'h4feefc3e7730;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[196] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[197] = 80'hd3f5a6c1574e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[197] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[198] = 80'hb6364f27da3b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[198] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[199] = 80'hdf1f0128cbbd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[199] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[200] = 80'h9cd060e84aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[200] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[201] = 80'h8373ac34c47f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[201] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[202] = 80'h1e386f8b863d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[202] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[203] = 80'h5ba2afce95f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[203] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[204] = 80'h4e2599a1897a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[204] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[205] = 80'hf5479d3b77c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[205] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[206] = 80'habbe127976b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[206] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[207] = 80'hda3b98564520;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[207] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[208] = 80'h5ac0acc44533;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[208] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[209] = 80'hddd77ea80899;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[209] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[210] = 80'h5ab30dbacc5d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[210] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[211] = 80'h342220f18625;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[211] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[212] = 80'h2a04827b867b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[212] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[213] = 80'h541f28ab2585;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[213] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[214] = 80'h283b331b6fc3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[214] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[215] = 80'h6f3ac91b9a16;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[215] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[216] = 80'h41fd7e0e3811;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[216] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[217] = 80'h58966af35810;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[217] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[218] = 80'he9cafeeb8643;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[218] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[219] = 80'hb3e98f6adfb5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[219] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[220] = 80'h739e76de29f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[220] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[221] = 80'h2a304169ea35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[221] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[222] = 80'h8151be21591a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[222] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[223] = 80'h1225f462349c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[223] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[224] = 80'h2719c0ef3496;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[224] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[225] = 80'h54fb7f3c0cef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[225] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[226] = 80'hfef0454047a7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[226] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[227] = 80'hb4d08228d18c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[227] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[228] = 80'ha167559cde76;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[228] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[229] = 80'h93813f42c579;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[229] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[230] = 80'h8510d813599c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[230] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[231] = 80'hd983360209d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[231] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[232] = 80'h9b211b4fc467;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[232] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[233] = 80'h2330c01b4962;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[233] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[234] = 80'h844df8e1f63b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[234] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[235] = 80'hc041ca14cdca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[235] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[236] = 80'hdaae12e7d039;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[236] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[237] = 80'h7036cba3dc70;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[237] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[238] = 80'hf19f6d156eb4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[238] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[239] = 80'h89fcfce01525;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[239] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[240] = 80'h1fad9639ae38;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[240] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[241] = 80'h59882292a37d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[241] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[242] = 80'hd1c038664adc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[242] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[243] = 80'h50d6e9dd8cb9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[243] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[244] = 80'h68165950944c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[244] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[245] = 80'hb1b417cc4d0d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[245] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[246] = 80'h673c0c16111e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[246] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[247] = 80'h9282fc16753b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[247] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[248] = 80'h465552830d4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[248] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[249] = 80'ha237c12459ce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[249] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[250] = 80'h3fbff4f63ebe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[250] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[251] = 80'h83622bea46ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[251] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[252] = 80'hace489475745;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[252] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[253] = 80'h1b62f58d5c3b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[253] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[254] = 80'h3d317dd9a17e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[254] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[255] = 80'h9b4487a8ad15;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[255] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[256] = 80'h1eb8f0ced706;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[256] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[257] = 80'h23df27639b89;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[257] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[258] = 80'h9e02d67f2c49;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[258] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[259] = 80'h2f03370d25d5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[259] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[260] = 80'h23c475b331f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[260] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[261] = 80'h298cf5b269e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[261] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[262] = 80'he8d802a6eec6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[262] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[263] = 80'hb112320fcf2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[263] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[264] = 80'h1e8b12608817;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[264] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[265] = 80'h70b74d52680c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[265] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[266] = 80'h9385b9ebc706;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[266] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[267] = 80'hc5ddaac7946a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[267] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[268] = 80'hd71073217127;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[268] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[269] = 80'hd100d643c643;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[269] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[270] = 80'hf69ca57a9df0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[270] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[271] = 80'hff6881bbfec2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[271] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[272] = 80'hf2823e7062c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[272] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[273] = 80'h61e0198f5ae3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[273] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[274] = 80'h2693612b76f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[274] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[275] = 80'h9e4433b3d0ed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[275] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[276] = 80'h1aa909a924ce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[276] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[277] = 80'h529bf4b7234;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[277] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[278] = 80'h71c5876f6f41;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[278] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[279] = 80'h4840ebc670dd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[279] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[280] = 80'he8a44e161d3a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[280] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[281] = 80'h45616bb46ded;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[281] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[282] = 80'h52dcbdb0812e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[282] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[283] = 80'h74514d0e52f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[283] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[284] = 80'h95635f45a99d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[284] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[285] = 80'h7ec8277acb2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[285] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[286] = 80'hdf530f8507d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[286] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[287] = 80'h76c5dc4ff347;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[287] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[288] = 80'hda63394fdb26;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[288] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[289] = 80'hdf60cec8ddc2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[289] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[290] = 80'h777e53ca6502;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[290] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[291] = 80'hfa9ef6faf654;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[291] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[292] = 80'he2fa7ff677c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[292] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[293] = 80'h1a6d4480a388;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[293] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[294] = 80'habf14b53db5d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[294] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[295] = 80'hd9e701d3b5a1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[295] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[296] = 80'hecb4c08dbedf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[296] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[297] = 80'h59425a4d73e4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[297] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[298] = 80'h46d500a7b842;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[298] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[299] = 80'h246ba174baea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[299] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[300] = 80'he1fa257edda3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[300] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[301] = 80'h9170e9535830;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[301] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[302] = 80'hb0da854090a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[302] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[303] = 80'h7794a452c0cc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[303] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[304] = 80'h1bb10373944d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[304] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[305] = 80'h54211c3f4263;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[305] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[306] = 80'h83f85a06a68f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[306] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[307] = 80'h262df1f69e49;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[307] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[308] = 80'h7d107f8ef4a6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[308] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[309] = 80'he4475d1bbe07;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[309] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[310] = 80'hf14033c3de26;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[310] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[311] = 80'heedc1c4b985;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[311] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[312] = 80'h45ea918b6353;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[312] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[313] = 80'hb6e8b1059138;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[313] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[314] = 80'he2d1f729b709;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[314] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[315] = 80'h358b6eaed36;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[315] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[316] = 80'ha67e6c68258f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[316] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[317] = 80'h3aa9c27a9590;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[317] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[318] = 80'h25062337c847;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[318] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[319] = 80'h2d9d36fde26f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[319] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[320] = 80'ha2f4f66c6e72;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[320] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[321] = 80'hd3dbc263b79e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[321] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[322] = 80'haa26b833ca5a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[322] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[323] = 80'he533d3adc92a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[323] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[324] = 80'he7989fff15b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[324] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[325] = 80'h204cb109b684;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[325] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[326] = 80'h9c86a3258c1c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[326] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[327] = 80'h33ee6b8cd041;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[327] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[328] = 80'h35cdd2ebe7d4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[328] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[329] = 80'hfbe9f071ba55;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[329] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[330] = 80'hedbaf396f94d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[330] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[331] = 80'h8f00c6959630;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[331] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[332] = 80'h2f0b7d02f677;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[332] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[333] = 80'h84361e779b29;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[333] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[334] = 80'hf9555655c72e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[334] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[335] = 80'h63fdd2831f64;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[335] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[336] = 80'h44f84811196a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[336] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[337] = 80'hee6a7ad1f326;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[337] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[338] = 80'hbd9a0d551dbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[338] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[339] = 80'hd77b6743a6d7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[339] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[340] = 80'hd514be473ad0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[340] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[341] = 80'hcd8d292c9163;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[341] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[342] = 80'h9b96c0a157f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[342] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[343] = 80'h3990be6ca74b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[343] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[344] = 80'h878954834a39;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[344] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[345] = 80'h55f55f90aaf2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[345] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[346] = 80'h6528fb359720;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[346] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[347] = 80'hd2e32bd26d81;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[347] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[348] = 80'h6cfb0768eaf9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[348] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[349] = 80'hf605651cbda8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[349] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[350] = 80'h67afeb283b90;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[350] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[351] = 80'h36956d2c31fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[351] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[352] = 80'heeff5a03dcc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[352] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[353] = 80'h68f890ba7165;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[353] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[354] = 80'h859e9ee2a203;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[354] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[355] = 80'h28b1629a2cd1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[355] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[356] = 80'hf9e13f57f9cb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[356] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[357] = 80'heb3232486a6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[357] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[358] = 80'h812ef34dfa60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[358] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[359] = 80'h390057c5b93d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[359] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[360] = 80'h9ebf1ea8a8a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[360] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[361] = 80'h3511debe665;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[361] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[362] = 80'h49fc818617e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[362] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[363] = 80'h9d37264bcd9f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[363] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[364] = 80'h9a822da69611;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[364] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[365] = 80'h27b44ca01d38;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[365] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[366] = 80'hc0c5608917d4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[366] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[367] = 80'h81edee6be9a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[367] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[368] = 80'h337d2f6ee9f6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[368] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[369] = 80'h3b0f04ce077f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[369] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[370] = 80'hfde55ff6a820;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[370] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[371] = 80'hdc321bcbeb8f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[371] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[372] = 80'h1bc1c7ca7403;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[372] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[373] = 80'hb7a0d02f7f9a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[373] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[374] = 80'h1c64b4b87959;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[374] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[375] = 80'h1e90fcb13925;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[375] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[376] = 80'h5ad1dcebe9aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[376] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[377] = 80'h45621e9591fb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[377] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[378] = 80'h59145ef9f8d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[378] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[379] = 80'h5605b54371f8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[379] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[380] = 80'hb963e37953dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[380] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[381] = 80'hd878910fbeb3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[381] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[382] = 80'he8578a861c2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[382] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[383] = 80'h4ec64f6caae0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[383] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[384] = 80'h854ba79d2364;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[384] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[385] = 80'h2cdf40fd45c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[385] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[386] = 80'ha01eaa448072;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[386] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[387] = 80'hd0441435aef0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[387] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[388] = 80'h5d2a8b0aef36;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[388] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[389] = 80'h8074ba3f6a36;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[389] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[390] = 80'h53797badc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[390] = 80'h7fffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[391] = 80'h2ed7fd573cf7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[391] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[392] = 80'he5883e982b3c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[392] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[393] = 80'h53a2748e29f6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[393] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[394] = 80'h5ca1a2544aa9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[394] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[395] = 80'he3f9ded7caed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[395] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[396] = 80'ha3643184f60a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[396] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[397] = 80'h2852f1edb5fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[397] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[398] = 80'h3244642a522c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[398] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[399] = 80'h577ae1143ac3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[399] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[400] = 80'hd116b38ae558;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[400] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[401] = 80'hef6f5c21938c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[401] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[402] = 80'hc7ae9723534c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[402] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[403] = 80'h12ee7fec5c3e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[403] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[404] = 80'h8ceb8fe138f0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[404] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[405] = 80'hac6c00b6a8d2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[405] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[406] = 80'hb15acb7a407c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[406] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[407] = 80'hfe01162b7c3d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[407] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[408] = 80'h3ca520daccf9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[408] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[409] = 80'h1ddba06c2730;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[409] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[410] = 80'h8c25018e78c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[410] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[411] = 80'h294e58af58b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[411] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[412] = 80'h25431f6f1ca8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[412] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[413] = 80'hd4e0d35b1bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[413] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[414] = 80'h288f8de89002;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[414] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[415] = 80'hbbd2142468fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[415] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[416] = 80'h9285b15180ce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[416] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[417] = 80'h89d7c1092a1f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[417] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[418] = 80'hbc5113c19cfc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[418] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[419] = 80'hcb0ad767c3ff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[419] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[420] = 80'h64d3dedd3b11;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[420] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[421] = 80'h1e5eb38233fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[421] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[422] = 80'hd9b98809ae51;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[422] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[423] = 80'h5f3093fd17e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[423] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[424] = 80'h8f220f87bb88;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[424] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[425] = 80'h2effec1166ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[425] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[426] = 80'h8efae6f79380;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[426] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[427] = 80'h1e1735b714f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[427] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[428] = 80'h74b95b6a5e36;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[428] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[429] = 80'had17df6d5280;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[429] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[430] = 80'hd9cc5ca6a92a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[430] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[431] = 80'hbcc4cdb632c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[431] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[432] = 80'h78702dc7b992;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[432] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[433] = 80'h4c0ae5cc4065;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[433] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[434] = 80'h6d192447580c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[434] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[435] = 80'h4082eb1df830;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[435] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[436] = 80'h6789fbb57be3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[436] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[437] = 80'h271e20654263;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[437] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[438] = 80'h46c0f48c2876;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[438] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[439] = 80'hb0e588475012;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[439] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[440] = 80'hf3bd582ea928;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[440] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[441] = 80'h2138e3a06726;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[441] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[442] = 80'ha916c7e72f2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[442] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[443] = 80'hb731cb59fe72;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[443] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[444] = 80'habcdc1e96b29;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[444] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[445] = 80'h38bcc2b05d26;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[445] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[446] = 80'h13f98cd1dbbd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[446] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[447] = 80'he592927a0a89;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[447] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[448] = 80'h9470cfe0bd38;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[448] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[449] = 80'hab62ba7b123c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[449] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[450] = 80'hc9793372f335;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[450] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[451] = 80'h17c05008dfd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[451] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[452] = 80'h7938cdcbad6d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[452] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[453] = 80'h282455e8a649;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[453] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[454] = 80'hd4b10f962ebd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[454] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[455] = 80'hee2a158883b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[455] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[456] = 80'h906a9ad30087;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[456] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[457] = 80'h4282827d137;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[457] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[458] = 80'h585a643eec07;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[458] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[459] = 80'heb073e9ed5c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[459] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[460] = 80'h21b4376f56e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[460] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[461] = 80'hbd2b7e328666;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[461] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[462] = 80'hf6b6101e438d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[462] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[463] = 80'h908022cd936f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[463] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[464] = 80'h7511ee9fa2de;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[464] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[465] = 80'h374776fb63b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[465] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[466] = 80'hd65c8503efa5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[466] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[467] = 80'h9ad572e1b926;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[467] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[468] = 80'h9e796c3e4446;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[468] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[469] = 80'h81296115c65e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[469] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[470] = 80'h2ef37672dd00;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[470] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[471] = 80'h1be09a9632b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[471] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[472] = 80'ha0251ac3bdd7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[472] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[473] = 80'hfa7f865e62ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[473] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[474] = 80'h290b9b7a1e05;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[474] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[475] = 80'h7f8e37e50737;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[475] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[476] = 80'he96a1056fbe0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[476] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[477] = 80'h492b7df8136d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[477] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[478] = 80'hb391bb6cff61;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[478] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[479] = 80'hb82153980608;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[479] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[480] = 80'habcbdbe195e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[480] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[481] = 80'hfcefb0d3fb08;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[481] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[482] = 80'h789711b0a797;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[482] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[483] = 80'h5cf2068e30a7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[483] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[484] = 80'hd4dfd545d947;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[484] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[485] = 80'h4926b200a921;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[485] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[486] = 80'hc373a403d24b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[486] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[487] = 80'h7e109be15c54;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[487] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[488] = 80'hb79c76af4364;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[488] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[489] = 80'h42ad91b91308;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[489] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[490] = 80'h923c87528181;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[490] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[491] = 80'h6927aecffc09;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[491] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[492] = 80'hb0d09ccc302d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[492] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[493] = 80'ha4234997ebd8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[493] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[494] = 80'h1ed04fa1ec97;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[494] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[495] = 80'h9892ee4621b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[495] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[496] = 80'hcfc813360aaa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[496] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[497] = 80'h5e383a86df15;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[497] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[498] = 80'h975c188f1dbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[498] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[499] = 80'h5ae15f494a6f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[499] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[500] = 80'hba60c9b84434;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[500] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[501] = 80'hec5378e383d8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[501] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[502] = 80'hc6f584a0c437;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[502] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[503] = 80'h37b198167e84;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[503] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[504] = 80'hd5a720e74827;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[504] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[505] = 80'h2b27ae1774a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[505] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[506] = 80'hd7ccbf2c8a33;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[506] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[507] = 80'hd7821106381a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[507] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[508] = 80'h27abf231a4f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[508] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[509] = 80'hf6b0f88997b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[509] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[510] = 80'h8bf13cd9575c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[510] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[511] = 80'h3269043ae182;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[511] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[512] = 80'ha08b34cab3ff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[512] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[513] = 80'h35f72570ae87;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[513] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[514] = 80'hef37fd8baffb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[514] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[515] = 80'hcaff585f4b5f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[515] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[516] = 80'h76eee9f3d2c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[516] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[517] = 80'haf06beec59cb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[517] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[518] = 80'h82c90775e233;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[518] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[519] = 80'hfe0847448447;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[519] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[520] = 80'hf0cb1f28c22a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[520] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[521] = 80'h7079f2078cc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[521] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[522] = 80'h6abd25be785f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[522] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[523] = 80'hdfdfc2f15c4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[523] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[524] = 80'hc9d15a930997;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[524] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[525] = 80'ha894e1e563f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[525] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[526] = 80'ha964fe119d5f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[526] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[527] = 80'h9dafde935b53;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[527] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[528] = 80'he906f4b5764;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[528] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[529] = 80'h216048dbe8e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[529] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[530] = 80'hc08f3732c7eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[530] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[531] = 80'hb72142bca4aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[531] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[532] = 80'h67a2ce8a5e0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[532] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[533] = 80'h5819e54162b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[533] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[534] = 80'hf81fb7436abb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[534] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[535] = 80'h31d8f5200247;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[535] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[536] = 80'h607df517446f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[536] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[537] = 80'h9501b95b8eee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[537] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[538] = 80'h4ac80e1571f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[538] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[539] = 80'h397eabef6f73;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[539] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[540] = 80'h58330b72f740;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[540] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[541] = 80'hb091099c5208;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[541] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[542] = 80'h8c922af3d544;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[542] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[543] = 80'h1ef54a94a1aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[543] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[544] = 80'heafb610d3307;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[544] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[545] = 80'h8f6e4315ccf3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[545] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[546] = 80'hbe335ca6def9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[546] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[547] = 80'hee0d6e2944d0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[547] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[548] = 80'hf79f7b4fbc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[548] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[549] = 80'h16a4b9b11745;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[549] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[550] = 80'hb854815e349a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[550] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[551] = 80'h8264f4b38d53;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[551] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[552] = 80'h2b31497dfe4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[552] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[553] = 80'h3874850e3664;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[553] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[554] = 80'h1e03504fc71e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[554] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[555] = 80'hac17c1eed961;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[555] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[556] = 80'h8b4a08190ea6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[556] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[557] = 80'h1a089420fe6b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[557] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[558] = 80'hdb0519d32d54;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[558] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[559] = 80'hd606b6890ccf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[559] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[560] = 80'h3a30d200a52e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[560] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[561] = 80'he1d629596d55;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[561] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[562] = 80'h59f8bd5018fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[562] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[563] = 80'h18c7b4420188;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[563] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[564] = 80'h381e1bed184a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[564] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[565] = 80'hd4a5ae2c135b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[565] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[566] = 80'he97961ccdcd0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[566] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[567] = 80'h737a13e21630;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[567] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[568] = 80'h6576d31493a8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[568] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[569] = 80'h16d47d0405e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[569] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[570] = 80'h33d13d02eaa0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[570] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[571] = 80'hd7950dbecaa4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[571] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[572] = 80'h58f7de01221a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[572] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[573] = 80'hf297721ec69a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[573] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[574] = 80'hfa8073a2c40f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[574] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[575] = 80'h991dda905a7c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[575] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[576] = 80'hb81a5d03ce28;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[576] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[577] = 80'h793b9c78b761;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[577] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[578] = 80'h48d383e9db0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[578] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[579] = 80'h94a5e12a8d29;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[579] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[580] = 80'h57351e593cda;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[580] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[581] = 80'h87cf3b2441aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[581] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[582] = 80'hf43a10956f47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[582] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[583] = 80'hde3fb55a35c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[583] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[584] = 80'h8018c8ac27bd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[584] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[585] = 80'h5a5c46dda87a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[585] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[586] = 80'h3c0309aa8715;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[586] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[587] = 80'h68918363bb53;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[587] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[588] = 80'h1a50f7d56556;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[588] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[589] = 80'h4141bcc97dea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[589] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[590] = 80'h30b786d0937c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[590] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[591] = 80'h4a0defcfa63e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[591] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[592] = 80'h4fefa8a8325b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[592] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[593] = 80'h65be949c2999;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[593] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[594] = 80'he228f54db17f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[594] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[595] = 80'hded2a0f4626e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[595] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[596] = 80'h43be668ec635;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[596] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[597] = 80'h642c6fad96e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[597] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[598] = 80'h869bf468988e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[598] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[599] = 80'h423d784e463c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[599] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[600] = 80'h9e0d7122e5d0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[600] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[601] = 80'hbbf5f3f9a3d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[601] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[602] = 80'h4d41bb7e83d4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[602] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[603] = 80'h9fe21480bf2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[603] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[604] = 80'h2daa4544c73c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[604] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[605] = 80'hde9abc1ba70d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[605] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[606] = 80'h74b4b8faa3cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[606] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[607] = 80'h53ffaa95bde0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[607] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[608] = 80'h7626b2b6c686;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[608] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[609] = 80'h63c350b895ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[609] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[610] = 80'hf4023a42fb3d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[610] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[611] = 80'hd063b376df50;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[611] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[612] = 80'hef9c58730d40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[612] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[613] = 80'hb7f07d70beeb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[613] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[614] = 80'hc6e6e5c33fca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[614] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[615] = 80'h32388657a2c4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[615] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[616] = 80'h6714ee2ee494;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[616] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[617] = 80'h95e542ea9383;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[617] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[618] = 80'h6ee62d6a2974;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[618] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[619] = 80'h992d98d8c860;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[619] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[620] = 80'h9d01df2dd16f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[620] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[621] = 80'h529561ddc2c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[621] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[622] = 80'hed170481df56;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[622] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[623] = 80'h8053bfce2d39;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[623] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[624] = 80'h2b3565e41eba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[624] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[625] = 80'hd039014a8676;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[625] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[626] = 80'h8aead6f8e415;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[626] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[627] = 80'hbc559f92bfc8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[627] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[628] = 80'h9ef7759a4335;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[628] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[629] = 80'h36050c4a38da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[629] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[630] = 80'h3a029f298309;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[630] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[631] = 80'hc13120cb0493;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[631] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[632] = 80'h4a807d566fcc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[632] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[633] = 80'hf4264c62ed60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[633] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[634] = 80'h60c439a2621c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[634] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[635] = 80'h66b493e0fe24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[635] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[636] = 80'h9b6927b93f7d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[636] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[637] = 80'h704b7af77695;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[637] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[638] = 80'h40ab28bca25f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[638] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[639] = 80'hc17bb0702ae1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[639] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[640] = 80'hb0d05cb346d2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[640] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[641] = 80'hcb0be3f40df1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[641] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[642] = 80'hb40e6c1f67e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[642] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[643] = 80'hdd08373eb7e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[643] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[644] = 80'h321f38e6c645;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[644] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[645] = 80'h22f54ffa712;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[645] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[646] = 80'h175711491a12;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[646] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[647] = 80'h5c4334e83dbf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[647] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[648] = 80'h7401586b796c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[648] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[649] = 80'h1064da257814;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[649] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[650] = 80'h33aa97849759;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[650] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[651] = 80'hdd749f6d10f2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[651] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[652] = 80'h32ec91b393dd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[652] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[653] = 80'h14cc9cebd56f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[653] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[654] = 80'hfa1a640d3120;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[654] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[655] = 80'hf4e3f6a941f0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[655] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[656] = 80'hd00f18748035;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[656] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[657] = 80'h471f97f6e335;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[657] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[658] = 80'h25d72449c9e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[658] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[659] = 80'h54f6d49980a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[659] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[660] = 80'hd9a3a9015e31;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[660] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[661] = 80'h7ca54a31df80;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[661] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[662] = 80'h2727fd6cbcb5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[662] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[663] = 80'h8d849e8d0bd6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[663] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[664] = 80'hc7917e2857fc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[664] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[665] = 80'hc114d4bda130;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[665] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[666] = 80'hbe6a2e10c1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[666] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[667] = 80'hef3b11cfca80;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[667] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[668] = 80'hda6802e720b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[668] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[669] = 80'hb955999acc64;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[669] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[670] = 80'hdc76ebecea5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[670] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[671] = 80'h3d59e483ea45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[671] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[672] = 80'h8e98064d1c2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[672] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[673] = 80'h111c13b657b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[673] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[674] = 80'hef7d1553096c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[674] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[675] = 80'h91047a599dcf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[675] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[676] = 80'ha8423d3eddb2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[676] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[677] = 80'hcfd34e86e5f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[677] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[678] = 80'h75ebdb494049;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[678] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[679] = 80'h3b3640c4d206;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[679] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[680] = 80'hd119b635c7bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[680] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[681] = 80'h719073427062;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[681] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[682] = 80'h5d2633c1c0c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[682] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[683] = 80'h5ffe5556f980;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[683] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[684] = 80'h61e8d059e1f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[684] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[685] = 80'h203ef10ced3e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[685] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[686] = 80'h9eee630d6efc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[686] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[687] = 80'h6322298a3a7b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[687] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[688] = 80'hf40c4bfc22fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[688] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[689] = 80'hfa5c7b97f665;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[689] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[690] = 80'hef9dfeb948eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[690] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[691] = 80'h382de4729315;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[691] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[692] = 80'h45bb0fa48950;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[692] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[693] = 80'h2ab5c380b341;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[693] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[694] = 80'h9f6273d1e971;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[694] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[695] = 80'hbc88ff2fe271;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[695] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[696] = 80'hc345fbecc076;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[696] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[697] = 80'hb6b2b6a8914d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[697] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[698] = 80'h69611d6f9e84;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[698] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[699] = 80'hbb21e0ea60b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[699] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem[700] = 80'h247897856c97;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[1].u_tcam.mem_mask[700] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[1] = 80'hc76428a3ac18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[1] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[2] = 80'h6fa2b332a044;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[2] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[3] = 80'hdf160ea7e244;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[3] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[4] = 80'hbde8a5158a2b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[4] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[5] = 80'h1c7fcaa5772f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[5] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[6] = 80'h398bc2065413;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[6] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[7] = 80'hbf26a132d23e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[7] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[8] = 80'h2e5a52ddfb3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[8] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[9] = 80'hf9c4f448c4c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[9] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[10] = 80'h35e4dd182f90;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[10] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[11] = 80'h8513d0c50521;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[11] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[12] = 80'h35a66285b62e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[12] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[13] = 80'h4915d9de428f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[13] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[14] = 80'h3eff489073c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[14] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[15] = 80'hd00165db49c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[15] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[16] = 80'hc6e7d540048a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[16] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[17] = 80'hd2cf31221e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[17] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[18] = 80'h9cc2400c08bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[18] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[19] = 80'he84ab68b1a24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[19] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[20] = 80'hdc9c606e91ae;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[20] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[21] = 80'h4b8ee53f7660;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[21] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[22] = 80'ha6dc109cdbbd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[22] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[23] = 80'h2e5acd726cb2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[23] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[24] = 80'hbb30b2ecd487;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[24] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[25] = 80'h9aeec82f8fac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[25] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[26] = 80'hab83fe2b985c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[26] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[27] = 80'hca3daac02b2f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[27] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[28] = 80'h1a893b2ffa10;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[28] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[29] = 80'hcb1ab883d9ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[29] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[30] = 80'h6ddb0412e88d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[30] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[31] = 80'h25d034a677c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[31] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[32] = 80'h2ee63ce89af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[32] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[33] = 80'h1ab5a710d843;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[33] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[34] = 80'h97e8c062f084;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[34] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[35] = 80'h30a809743d4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[35] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[36] = 80'h22420da7f8f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[36] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[37] = 80'hafaf284ad3bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[37] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[38] = 80'h53bd4f0d7794;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[38] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[39] = 80'h5c0d39f2f061;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[39] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[40] = 80'h9419a7ce074a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[40] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[41] = 80'h52d45cc1e4a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[41] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[42] = 80'h9b30665b9971;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[42] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[43] = 80'h20d936f412c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[43] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[44] = 80'h8b889af41550;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[44] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[45] = 80'hf91ce85e797d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[45] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[46] = 80'h6e1dbd81191;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[46] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[47] = 80'h345e3c5f1365;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[47] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[48] = 80'h8dceefe91dc9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[48] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[49] = 80'hd47d2191ffed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[49] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[50] = 80'h7d341fbc821b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[50] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[51] = 80'h2e1c5d9ff7d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[51] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[52] = 80'hb7c667fd0324;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[52] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[53] = 80'h4933bf21a16c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[53] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[54] = 80'hf9724902347e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[54] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[55] = 80'haeb766b220db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[55] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[56] = 80'hdbbc2a3224ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[56] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[57] = 80'h365a679e8085;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[57] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[58] = 80'heeff7c2b7b33;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[58] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[59] = 80'h45bb6a31bb68;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[59] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[60] = 80'h1a81b1c43f91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[60] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[61] = 80'h1de0ad29184a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[61] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[62] = 80'h4eb9229cd415;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[62] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[63] = 80'h75c39cfd15db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[63] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[64] = 80'hbd7d9ddf726;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[64] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[65] = 80'h788ece7eed43;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[65] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[66] = 80'h689790000fff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[66] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[67] = 80'h30fca31cf96b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[67] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[68] = 80'h358975cc2823;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[68] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[69] = 80'h6b1cd921c79d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[69] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[70] = 80'h549a31ff63b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[70] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[71] = 80'h310dee607220;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[71] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[72] = 80'haf90fc2fb606;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[72] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[73] = 80'hdb655000d3a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[73] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[74] = 80'h8bf35344ab45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[74] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[75] = 80'h2d8a38190b20;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[75] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[76] = 80'h263f7f66582;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[76] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[77] = 80'h4dfc2ba4768d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[77] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[78] = 80'h849983bfbe7a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[78] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[79] = 80'h1efcb2f4dd4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[79] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[80] = 80'h61e5a9de4569;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[80] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[81] = 80'h770c1c4bd3a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[81] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[82] = 80'h500562660aff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[82] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[83] = 80'ha72a189143e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[83] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[84] = 80'h51a64abf0e09;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[84] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[85] = 80'h1f5700abe928;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[85] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[86] = 80'h512e72fad6a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[86] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[87] = 80'h5f3a530396cf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[87] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[88] = 80'h748487400445;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[88] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[89] = 80'h87719fb3f864;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[89] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[90] = 80'he88c8f60061d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[90] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[91] = 80'h9f6cc5f93019;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[91] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[92] = 80'hfa9df2c0fa11;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[92] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[93] = 80'h3e5de237f4f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[93] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[94] = 80'h1220e6f8b9fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[94] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[95] = 80'hceb0c2f94c3c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[95] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[96] = 80'h1845b8356ded;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[96] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[97] = 80'hcb7d6f052ed9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[97] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[98] = 80'ha1d827523dc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[98] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[99] = 80'hcaf8264a3ea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[99] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[100] = 80'h38ead3f12916;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[100] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[101] = 80'h13d2ee37c448;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[101] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[102] = 80'h3c2fe7d9f34c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[102] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[103] = 80'h3c1db8626079;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[103] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[104] = 80'h865b861ca607;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[104] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[105] = 80'h794600c6d0f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[105] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[106] = 80'he00c57f6e0b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[106] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[107] = 80'he29db65e8903;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[107] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[108] = 80'h8e261e6170f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[108] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[109] = 80'h66939b10ec73;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[109] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[110] = 80'h70c2e9c3c8eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[110] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[111] = 80'h45c66be84cf4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[111] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[112] = 80'h232cef211d0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[112] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[113] = 80'h80542dda5aa2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[113] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[114] = 80'h474effbc30dd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[114] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[115] = 80'he4cebd5c6fa4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[115] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[116] = 80'haf6a54830375;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[116] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[117] = 80'h8ef028be44c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[117] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[118] = 80'h5fdca8436bf4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[118] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[119] = 80'h6e7e1c15bd08;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[119] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[120] = 80'h134c1f65fd66;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[120] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[121] = 80'hcea87493679f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[121] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[122] = 80'hceb7bc309c1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[122] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[123] = 80'h61a6f8771878;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[123] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[124] = 80'hcedef6a567fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[124] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[125] = 80'h2e32a08622cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[125] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[126] = 80'h5356e16b8fd7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[126] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[127] = 80'hfd605bd942c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[127] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[128] = 80'hd5f103f449;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[128] = 80'hffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[129] = 80'h5f57f4362b22;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[129] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[130] = 80'h2e67f284f871;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[130] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[131] = 80'hecd79dcadc01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[131] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[132] = 80'he00525c7b0f8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[132] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[133] = 80'hb3cf483e6c80;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[133] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[134] = 80'h77eb26f31bbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[134] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[135] = 80'h8b676c49d915;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[135] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[136] = 80'ha2822acbd35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[136] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[137] = 80'h3a257929df1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[137] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[138] = 80'he9b0e1c40a18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[138] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[139] = 80'h3f10a0b32f42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[139] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[140] = 80'hf8a042a8b1d1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[140] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[141] = 80'hc010041f98fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[141] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[142] = 80'h6f5155d6bf2a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[142] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[143] = 80'h6174e0aee88e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[143] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[144] = 80'hd8f296505931;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[144] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[145] = 80'he512e3c64789;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[145] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[146] = 80'h373e0b9976b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[146] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[147] = 80'h3e7dacda18b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[147] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[148] = 80'h964ddbc00a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[148] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[149] = 80'h54781b947c65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[149] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[150] = 80'h4e476ae23070;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[150] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[151] = 80'h965a202c5dd1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[151] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[152] = 80'h6eeef25e5a0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[152] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[153] = 80'hbd9be825e53c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[153] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[154] = 80'h5a0d2b0e2652;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[154] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[155] = 80'hf02c2960a78f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[155] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[156] = 80'h43801573ed5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[156] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[157] = 80'h34d1a3628645;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[157] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[158] = 80'h476d2c7ebc16;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[158] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[159] = 80'ha17de6c9b9c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[159] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[160] = 80'h2e3b2da7cb0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[160] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[161] = 80'h618fe75b3a00;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[161] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[162] = 80'h7868e9b929a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[162] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[163] = 80'hcbe5e4137d1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[163] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[164] = 80'h6771e8c490b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[164] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[165] = 80'h7be9cc15dbad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[165] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[166] = 80'h8c89b097b14c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[166] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[167] = 80'hf2124342ae18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[167] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[168] = 80'h330261ba3670;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[168] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[169] = 80'h42c4edb6d896;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[169] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[170] = 80'h23a570bc32da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[170] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[171] = 80'hdb4f2973fc73;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[171] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[172] = 80'h4c40d88318b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[172] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[173] = 80'h1273739101e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[173] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[174] = 80'h9c2ebac8770d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[174] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[175] = 80'haaeaffde1744;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[175] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[176] = 80'h67b1d0406ac4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[176] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[177] = 80'h602be7c25423;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[177] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[178] = 80'h7bd2374d89da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[178] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[179] = 80'h484efbf68ee5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[179] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[180] = 80'h8c2970d5df55;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[180] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[181] = 80'haec65cebfe7b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[181] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[182] = 80'h94dfc4cad63a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[182] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[183] = 80'h16398c9c5329;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[183] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[184] = 80'hc1d9c5b84501;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[184] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[185] = 80'hd1ad3332662b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[185] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[186] = 80'hb91d094ca5fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[186] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[187] = 80'h66807169ce5b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[187] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[188] = 80'h6ef096e4f564;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[188] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[189] = 80'h328864e675f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[189] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[190] = 80'h7dae2b0e1b45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[190] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[191] = 80'hbcb94b47b6e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[191] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[192] = 80'h969630df4be5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[192] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[193] = 80'h8fa1021a531a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[193] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[194] = 80'h872d61d5debf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[194] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[195] = 80'h991610788933;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[195] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[196] = 80'habf899e0a35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[196] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[197] = 80'h9a50b37b4c4e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[197] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[198] = 80'ha57859f9c477;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[198] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[199] = 80'h79cd60c49c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[199] = 80'h7fffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[200] = 80'h116a5a1abd7d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[200] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[201] = 80'hc21fd0b46818;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[201] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[202] = 80'hcb7c1d8cfffa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[202] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[203] = 80'h5da2668e789f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[203] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[204] = 80'ha975554d1660;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[204] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[205] = 80'hf527f8412a24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[205] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[206] = 80'h6e7cabe12a47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[206] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[207] = 80'hecce1c4cd86e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[207] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[208] = 80'h72d3d3fcd72b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[208] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[209] = 80'h839e1fb55d44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[209] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[210] = 80'h478398e0b9ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[210] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[211] = 80'h8530d50e759f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[211] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[212] = 80'h11f968361ebd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[212] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[213] = 80'h8ce994cc083f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[213] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[214] = 80'h2c23f84988ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[214] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[215] = 80'h9760938f25c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[215] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[216] = 80'h274efbfa8211;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[216] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[217] = 80'h694132b93ba3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[217] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[218] = 80'h682f3056401;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[218] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[219] = 80'hd1c36a785d4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[219] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[220] = 80'h4ae9b6d2ef4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[220] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[221] = 80'hc9c32ab41eeb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[221] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[222] = 80'hcbc076ebe28e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[222] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[223] = 80'hfbda31fd76c0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[223] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[224] = 80'h9a099a151b35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[224] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[225] = 80'h54a1681b3ffb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[225] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[226] = 80'hf0cf8f9ee272;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[226] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[227] = 80'h3f535b44d28a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[227] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[228] = 80'h7ae44fa333c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[228] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[229] = 80'hb665ce7f735a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[229] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[230] = 80'h626c7ae8774d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[230] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[231] = 80'hf3cddb51d392;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[231] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[232] = 80'h944a75a8319c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[232] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[233] = 80'heaacb9890fae;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[233] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[234] = 80'h46f6540ec7f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[234] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[235] = 80'hc6088fc1bd3d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[235] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[236] = 80'h5e0b61c56031;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[236] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[237] = 80'h27b4c51c3bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[237] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[238] = 80'hbe4d82d7e60e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[238] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[239] = 80'h7eef6a0932c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[239] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[240] = 80'h564f40cb3bc6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[240] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[241] = 80'h49ba0e14ede1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[241] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[242] = 80'hffa1385e8e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[242] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[243] = 80'hc2a6a6c5875c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[243] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[244] = 80'h46ed88992ff9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[244] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[245] = 80'h7bd52c488741;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[245] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[246] = 80'hdd037b320186;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[246] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[247] = 80'hbc45bae8ac0a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[247] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[248] = 80'h5b06c7e96f30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[248] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[249] = 80'hd4ddc557a673;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[249] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[250] = 80'h53ec21af6aa7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[250] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[251] = 80'h17ac57f88e87;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[251] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[252] = 80'ha4100e4032cc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[252] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[253] = 80'h140fa51dda60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[253] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[254] = 80'hba76b63b04af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[254] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[255] = 80'h7bf30212d42d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[255] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[256] = 80'h389a856d0929;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[256] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[257] = 80'h971def77bfa0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[257] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[258] = 80'h7fea6ca2dda9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[258] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[259] = 80'h6cc87b7163e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[259] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[260] = 80'h652f37432033;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[260] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[261] = 80'h94ca0afeaf40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[261] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[262] = 80'haa6075a82cfd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[262] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[263] = 80'he393132fbd4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[263] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[264] = 80'h8617fb8769a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[264] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[265] = 80'hd45704f554fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[265] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[266] = 80'h83aeac67707;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[266] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[267] = 80'had11dd592c9a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[267] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[268] = 80'h199fcd09ed28;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[268] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[269] = 80'h306fc67d4fd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[269] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[270] = 80'hded308236673;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[270] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[271] = 80'h6bb4f3981543;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[271] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[272] = 80'h28d774fa8bab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[272] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[273] = 80'h5f39e126fa40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[273] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[274] = 80'h4ec1930dd830;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[274] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[275] = 80'h2eabafa47444;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[275] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[276] = 80'hf2c4354979b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[276] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[277] = 80'h4375ff2839ff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[277] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[278] = 80'h831847d750e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[278] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[279] = 80'h6d4ff70a7fc3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[279] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[280] = 80'h67633ad96690;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[280] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[281] = 80'h58b1bb7ab35b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[281] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[282] = 80'h378d65b1297a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[282] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[283] = 80'h8ab24a720a34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[283] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[284] = 80'h9b617faf808a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[284] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[285] = 80'h2b5be33345f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[285] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[286] = 80'h80b069925240;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[286] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[287] = 80'h64819ae5ce38;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[287] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[288] = 80'hc8a2886319ad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[288] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[289] = 80'hbba80680cd74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[289] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[290] = 80'hc624c1780420;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[290] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[291] = 80'hdf4dc19f8a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[291] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[292] = 80'hbf4fc4c5109d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[292] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[293] = 80'h230e53a6e40d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[293] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[294] = 80'h6a8845704812;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[294] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[295] = 80'hd02d7e61c3ff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[295] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[296] = 80'h42d9ad4b7cb5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[296] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[297] = 80'h6620c43e40cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[297] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[298] = 80'h572b2a5075a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[298] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[299] = 80'hbc0a3cd8632;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[299] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[300] = 80'h318840f45c23;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[300] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[301] = 80'h7ec0b9f2df84;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[301] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[302] = 80'h708eaeea371;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[302] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[303] = 80'h29e3e9901c1f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[303] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[304] = 80'hf4f0fb40376f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[304] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[305] = 80'h7de8c27c7bf8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[305] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[306] = 80'h722214538bb3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[306] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[307] = 80'hb35284a2e8f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[307] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[308] = 80'hc1e963dc4088;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[308] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[309] = 80'h50d5503770e6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[309] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[310] = 80'hb63951662a30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[310] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[311] = 80'h7eddea567619;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[311] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[312] = 80'h4eab0a109e8f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[312] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[313] = 80'he549f26a551a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[313] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[314] = 80'h161e12d7d5f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[314] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[315] = 80'h2fb8691cf03d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[315] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[316] = 80'h6d0dd414bd88;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[316] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[317] = 80'hd47f0cfd8269;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[317] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[318] = 80'he7fe58f76aac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[318] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[319] = 80'hcddb5437e4b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[319] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[320] = 80'h58ac2d7d65c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[320] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[321] = 80'he81d8eb85034;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[321] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[322] = 80'ha6fb99d69d1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[322] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[323] = 80'h85db0f2ad52e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[323] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[324] = 80'hba447f49c0b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[324] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[325] = 80'h99d3496acd35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[325] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[326] = 80'h40e7e1b07303;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[326] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[327] = 80'h55f948ebe91d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[327] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[328] = 80'h392c0459ce02;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[328] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[329] = 80'h7e3d419f5d34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[329] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[330] = 80'he74efb58eaa7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[330] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[331] = 80'hf83f581e4482;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[331] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[332] = 80'h9cce1dfeef14;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[332] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[333] = 80'h4b70936e9f64;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[333] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[334] = 80'h8f60bf446783;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[334] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[335] = 80'h93a9046448e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[335] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[336] = 80'h6e3ce4ac6730;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[336] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[337] = 80'h84de22fbc40a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[337] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[338] = 80'h2d98732c0914;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[338] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[339] = 80'h588e0584287c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[339] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[340] = 80'h8f50e0497e89;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[340] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[341] = 80'hb0e119fb2555;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[341] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[342] = 80'h4cd3c2cde21a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[342] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[343] = 80'hda342cb3beee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[343] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[344] = 80'h9f7fc5e6a042;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[344] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[345] = 80'hcc5300c82669;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[345] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[346] = 80'h6a1ec386bf00;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[346] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[347] = 80'h2317e8d90545;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[347] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[348] = 80'h8d4fe98625cf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[348] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[349] = 80'h60665e2c19e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[349] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[350] = 80'h596674fbbfb1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[350] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[351] = 80'h5c7688d8aad5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[351] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[352] = 80'h99c3cb202d30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[352] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[353] = 80'ha86ac83a7681;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[353] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[354] = 80'hf9f330aaf7e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[354] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[355] = 80'h3c3dcdb988e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[355] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[356] = 80'h82440e73e0a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[356] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[357] = 80'hdeb63d376bdd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[357] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[358] = 80'h3f13c6d986da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[358] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[359] = 80'h959a11161a8a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[359] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[360] = 80'h4fc4b9709a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[360] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[361] = 80'h603260a4fa8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[361] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[362] = 80'h317642426d30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[362] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[363] = 80'h93eea5159da0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[363] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[364] = 80'ha6a6c5effbb8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[364] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[365] = 80'h9a556fc0f1e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[365] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[366] = 80'hca8bfde422b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[366] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[367] = 80'h6b3d4da4a0e4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[367] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[368] = 80'hb8725432eee0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[368] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[369] = 80'h2a5f4d97572c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[369] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[370] = 80'h3f4b2f37c91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[370] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[371] = 80'h6d012a56f306;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[371] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[372] = 80'hf39c18ff7423;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[372] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[373] = 80'h64fe54c3d020;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[373] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[374] = 80'h5941386df853;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[374] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[375] = 80'hfd5081a7023d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[375] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[376] = 80'h59d252677e44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[376] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[377] = 80'hb1ef710456c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[377] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[378] = 80'h8a3b29afa55f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[378] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[379] = 80'ha8f4af7c920a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[379] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[380] = 80'h9b5b556528f0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[380] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[381] = 80'h8d75c4ce6384;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[381] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[382] = 80'h644e172a4d39;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[382] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[383] = 80'h4e2c31c4e9bf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[383] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[384] = 80'hfb16e104670e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[384] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[385] = 80'hedda66338267;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[385] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[386] = 80'h28c12a16f1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[386] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[387] = 80'hff84824ad314;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[387] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[388] = 80'hbe7756aeeab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[388] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[389] = 80'h7e61e055303f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[389] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[390] = 80'haac7193a22af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[390] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[391] = 80'h565f0106873e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[391] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[392] = 80'h75032e61802d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[392] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[393] = 80'hf2f7c9dbbf6e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[393] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[394] = 80'hc616b82074dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[394] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[395] = 80'h9b90c73a26b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[395] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[396] = 80'hf1aad48501e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[396] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[397] = 80'hb50e5a5b2331;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[397] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[398] = 80'h536e70ff511;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[398] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[399] = 80'h500f137223d6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[399] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[400] = 80'h2791051b62a6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[400] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[401] = 80'hc4eb2c045df0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[401] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[402] = 80'ha4ad1b4e4c65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[402] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[403] = 80'h5dcd203c62ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[403] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[404] = 80'hbd2053fe1aa1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[404] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[405] = 80'hdd873733eebd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[405] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[406] = 80'hd5cc8944cc44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[406] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[407] = 80'hdf75e34c1d60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[407] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[408] = 80'h69516c90e02b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[408] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[409] = 80'hba7434218648;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[409] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[410] = 80'h75995e082cc9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[410] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[411] = 80'h8f8a0618c492;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[411] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[412] = 80'h85652adefb50;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[412] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[413] = 80'h84e3bbb346a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[413] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[414] = 80'hce288545ff5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[414] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[415] = 80'hf34840529bc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[415] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[416] = 80'h93b680734ca8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[416] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[417] = 80'h6d3e5930bf31;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[417] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[418] = 80'h4c6bb4e13dd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[418] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[419] = 80'hc17e7cae146d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[419] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[420] = 80'h3a01e234f448;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[420] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[421] = 80'h1f6089a70d31;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[421] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[422] = 80'he9910acedf01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[422] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[423] = 80'h92c1be63a45c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[423] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[424] = 80'h77250b5545e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[424] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[425] = 80'h41875a4af1b4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[425] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[426] = 80'h1f7188b8f195;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[426] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[427] = 80'he7043697f5e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[427] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[428] = 80'hccb0a5325cbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[428] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[429] = 80'hf77c99d0ae10;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[429] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[430] = 80'h51c66267cec7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[430] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[431] = 80'ha3eb7b517f7d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[431] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[432] = 80'h5e4b84a9a324;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[432] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[433] = 80'h263366d9a934;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[433] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[434] = 80'h35cd167e2bad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[434] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[435] = 80'hb2c3bbf8fba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[435] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[436] = 80'h8f19a66976c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[436] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[437] = 80'he0b42c35622b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[437] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[438] = 80'hdca9a6f1782c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[438] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[439] = 80'h9a1541c274a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[439] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[440] = 80'h44768a38b95d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[440] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[441] = 80'h38f48a68b142;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[441] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[442] = 80'h9759c188b4fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[442] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[443] = 80'ha08c0f3399b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[443] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[444] = 80'h820dea118ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[444] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[445] = 80'h786f4fec3569;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[445] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[446] = 80'h35502a9bf339;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[446] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[447] = 80'hede032f81911;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[447] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[448] = 80'h5d2da41d57;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[448] = 80'h7fffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[449] = 80'h1d551e45233a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[449] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[450] = 80'h1232e7e21619;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[450] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[451] = 80'h9656bf8e0b9d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[451] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[452] = 80'h282df63c9a42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[452] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[453] = 80'hfb8cfa3efc1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[453] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[454] = 80'he202a5e04142;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[454] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[455] = 80'hce14bd93ed55;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[455] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[456] = 80'hb29b6b75332;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[456] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[457] = 80'ha560cfe7acfc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[457] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[458] = 80'h99c7f0448e01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[458] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[459] = 80'h1dc007e9c85a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[459] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[460] = 80'hd5bbfcebded1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[460] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[461] = 80'h7a59ce859cc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[461] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[462] = 80'h4ea8c5b70bda;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[462] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[463] = 80'h52f1807fc08a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[463] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[464] = 80'h206171d9529a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[464] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[465] = 80'h498a7ea9d6a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[465] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[466] = 80'h68b1d8990008;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[466] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[467] = 80'hdfdd7f5c6649;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[467] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[468] = 80'h423c83f43d47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[468] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[469] = 80'h71daa74440c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[469] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[470] = 80'h6b7caeb2cb69;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[470] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[471] = 80'h9301716b199f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[471] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[472] = 80'hf30c2c261355;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[472] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[473] = 80'he1037b5789b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[473] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[474] = 80'h4ac85c163c30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[474] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[475] = 80'hbd2e17a3bd71;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[475] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[476] = 80'h8cfbaac12a25;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[476] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[477] = 80'he07f86b355a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[477] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[478] = 80'he24b3b5f435d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[478] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[479] = 80'hc6100a3221e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[479] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[480] = 80'hd601e9e5d6ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[480] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[481] = 80'ha2ee82f9007b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[481] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[482] = 80'hb4baf8944204;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[482] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[483] = 80'h78c5ee1f506d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[483] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[484] = 80'h94176a64d950;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[484] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[485] = 80'hbdc7edf2bed3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[485] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[486] = 80'hf6141087125a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[486] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[487] = 80'h4d8a6c4bb175;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[487] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[488] = 80'hd702b7ff755e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[488] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[489] = 80'h17ad459c4491;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[489] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[490] = 80'hbecd69de0af5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[490] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[491] = 80'h6db83a09cb40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[491] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[492] = 80'hc15a3192c54e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[492] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[493] = 80'h372729de79a7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[493] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[494] = 80'hb7d5a573112e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[494] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[495] = 80'he7598a8d64ef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[495] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[496] = 80'h4d77a8f186e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[496] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[497] = 80'hb3a7e8c62438;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[497] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[498] = 80'h5e628e40bad8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[498] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[499] = 80'h2c6ae9566a81;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[499] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[500] = 80'h7c8088a4d780;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[500] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[501] = 80'h449da718991b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[501] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[502] = 80'heb14915c851e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[502] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[503] = 80'h3527b3d245b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[503] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[504] = 80'h85d7cc131a8a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[504] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[505] = 80'hb448dcc734b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[505] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[506] = 80'h463282aaf56;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[506] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[507] = 80'he6f6fe35b667;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[507] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[508] = 80'h80c258b15826;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[508] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[509] = 80'hfaac4f7283f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[509] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[510] = 80'ha03cce697a88;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[510] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[511] = 80'hdf03c7e186d0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[511] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[512] = 80'hc301b2ddb491;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[512] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[513] = 80'h5a553a6d946;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[513] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[514] = 80'hec81a0ecf565;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[514] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[515] = 80'h25b7ba6c7a22;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[515] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[516] = 80'hff62f77af68e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[516] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[517] = 80'h90696c0e7c49;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[517] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[518] = 80'hdb542752b51b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[518] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[519] = 80'h5c669d7e5719;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[519] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[520] = 80'h7869b90d6d6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[520] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[521] = 80'h6ab3f4028bc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[521] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[522] = 80'hfaf254c81784;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[522] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[523] = 80'he91e80ddf2b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[523] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[524] = 80'h12ec8002dccf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[524] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[525] = 80'h1fb66119b301;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[525] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[526] = 80'h35cfa56dca6a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[526] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[527] = 80'h257f17287640;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[527] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[528] = 80'he24b719e5fd5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[528] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[529] = 80'h1b6de98d63bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[529] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[530] = 80'hc7396a1e1d0b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[530] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[531] = 80'h7fb43ae9cd4b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[531] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[532] = 80'ha389a8825008;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[532] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[533] = 80'h62002cc089d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[533] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[534] = 80'ha2fc3e097fd8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[534] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[535] = 80'h93938f2e7bb6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[535] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[536] = 80'h4c0878c8f3c9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[536] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[537] = 80'h6dad4681d74b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[537] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[538] = 80'h90d849afd440;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[538] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[539] = 80'h99cea5c192b2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[539] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[540] = 80'h439a63924ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[540] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[541] = 80'h22efe4c3db4e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[541] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[542] = 80'h935f8ae1eaca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[542] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[543] = 80'h980ce89cb3ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[543] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[544] = 80'hb2b1d54e6143;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[544] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[545] = 80'h985262ca09c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[545] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[546] = 80'h1b5370c23148;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[546] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[547] = 80'hfa6e44897737;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[547] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[548] = 80'hedc347b5f551;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[548] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[549] = 80'hbbafbcb86844;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[549] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[550] = 80'h7fb9ba95cb59;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[550] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[551] = 80'hbe931b35ee21;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[551] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[552] = 80'h39f56d709e34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[552] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[553] = 80'h4e9dfa08200a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[553] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[554] = 80'h820c31b21a45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[554] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[555] = 80'h5c7809f7005;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[555] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[556] = 80'h3aca0c094cca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[556] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[557] = 80'h745ae42f60b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[557] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[558] = 80'h9ab1034e7c6e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[558] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[559] = 80'h8b03e00b02c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[559] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[560] = 80'h291393c268aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[560] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[561] = 80'h4f5dda910b46;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[561] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[562] = 80'hd702572b740;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[562] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[563] = 80'h82eb751a50eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[563] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[564] = 80'h69f1bf212be5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[564] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[565] = 80'h692f8eeae2e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[565] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[566] = 80'h19a683169415;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[566] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[567] = 80'h93bac3e6e685;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[567] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[568] = 80'h4993bee769ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[568] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[569] = 80'hcd7fb4cb6753;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[569] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[570] = 80'h240e7a3c36d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[570] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[571] = 80'hdee7cb29be85;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[571] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[572] = 80'h992597565e42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[572] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[573] = 80'h5cf48819c736;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[573] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[574] = 80'h47abe210da7f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[574] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[575] = 80'hf93a1757baa0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[575] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[576] = 80'h7c1ceb4afc56;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[576] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[577] = 80'haf7d256d7cc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[577] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[578] = 80'h56f4eacb32c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[578] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[579] = 80'hb0d1add53e47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[579] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[580] = 80'hd2755cc4bd17;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[580] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[581] = 80'ha6985589f9f2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[581] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[582] = 80'hc617a79d7ece;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[582] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[583] = 80'hce74602fffba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[583] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[584] = 80'hf924b4b96d61;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[584] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[585] = 80'h8c0b6b9901dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[585] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[586] = 80'hf68af87708bf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[586] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[587] = 80'h74fa5f30fe3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[587] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[588] = 80'h4db8a921b1d2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[588] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[589] = 80'h18a72f979e24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[589] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[590] = 80'h595e18260e26;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[590] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[591] = 80'haad2d483e822;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[591] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[592] = 80'h343913fad305;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[592] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[593] = 80'hb3d2b6c10e97;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[593] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[594] = 80'h5b359f4f70b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[594] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[595] = 80'h910fdf65238e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[595] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[596] = 80'h858d2a03d342;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[596] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[597] = 80'h60c0b6079327;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[597] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[598] = 80'hac7bf03559d7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[598] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[599] = 80'h9ad2390bbe32;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[599] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[600] = 80'hfa4f7ce06718;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[600] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[601] = 80'hd16fe65ec39f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[601] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[602] = 80'h2d99e55053a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[602] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[603] = 80'h5159029f3697;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[603] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[604] = 80'hb4b0447b5549;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[604] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[605] = 80'h377b752a37b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[605] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[606] = 80'h220bb11437f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[606] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[607] = 80'habd69fb1204e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[607] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[608] = 80'heb47988d0d8b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[608] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[609] = 80'hca9cc767edce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[609] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[610] = 80'h3b6f42cbe0a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[610] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[611] = 80'h1dd3fa287076;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[611] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[612] = 80'h9628912dbff2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[612] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[613] = 80'h89a7951bea35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[613] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[614] = 80'hc7b2ff90ab75;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[614] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[615] = 80'h7ec37d3f35d1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[615] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[616] = 80'h486d45350ba4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[616] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[617] = 80'hf7c78a4aeffd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[617] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[618] = 80'hea7f3c4470a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[618] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[619] = 80'h95398bca46db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[619] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[620] = 80'h2a21d269ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[620] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[621] = 80'h5ff142432afa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[621] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[622] = 80'h8d346fc65e2b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[622] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[623] = 80'h1a6584f50556;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[623] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[624] = 80'h8386da1029f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[624] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[625] = 80'hdb56c981ece6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[625] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[626] = 80'hcfe8af38f522;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[626] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[627] = 80'h8e919d8a745b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[627] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[628] = 80'h543818958c78;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[628] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[629] = 80'ha8b931f97188;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[629] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[630] = 80'h7dee0d849922;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[630] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[631] = 80'h1017ca8a2953;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[631] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[632] = 80'h7ed9cae24403;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[632] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[633] = 80'hea187ed4d55a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[633] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[634] = 80'h2e76e28270f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[634] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[635] = 80'hf1980343333f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[635] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[636] = 80'h8de1c963c062;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[636] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[637] = 80'h3fd86ea44501;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[637] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[638] = 80'hdc791a00bf2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[638] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[639] = 80'h76fd772b3105;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[639] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[640] = 80'h9137a6d429b2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[640] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[641] = 80'h49d4cbef7ccc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[641] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[642] = 80'h8051f12b529f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[642] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[643] = 80'h8d6aa657a5e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[643] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[644] = 80'h44bafb829ee6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[644] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[645] = 80'he55061ccc7b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[645] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[646] = 80'hd75970bd3bb0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[646] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[647] = 80'h4811729ba385;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[647] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[648] = 80'hc0501fd955df;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[648] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[649] = 80'h659c29b06d69;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[649] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[650] = 80'h6aec373261a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[650] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[651] = 80'hc25cd90f5dab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[651] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[652] = 80'hcee3230bfef6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[652] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[653] = 80'h7bde198a992f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[653] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[654] = 80'h7cd4d9587ccb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[654] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[655] = 80'h5cee7e94dd42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[655] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[656] = 80'hc7f2c96b613;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[656] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[657] = 80'hf2de9d0bdde4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[657] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[658] = 80'hb80342294761;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[658] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[659] = 80'hef05f9051dde;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[659] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[660] = 80'h89d9864b0f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[660] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[661] = 80'hf84ebc6b5933;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[661] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[662] = 80'h99c7ebd6ef11;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[662] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[663] = 80'ha5cfc726453c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[663] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[664] = 80'h8e33ccc43905;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[664] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[665] = 80'h61dbc393f8b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[665] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[666] = 80'hb5776eb8e40c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[666] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[667] = 80'hc56f02fbb8af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[667] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[668] = 80'hf06ac89a6e2e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[668] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[669] = 80'h4d46ea5704c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[669] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[670] = 80'h18a0d2ab536;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[670] = 80'h1ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[671] = 80'hde24ea9c8559;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[671] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[672] = 80'h117c2dcb8a3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[672] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[673] = 80'h42c5800a198;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[673] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[674] = 80'hc866641162c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[674] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[675] = 80'hc59ce2a178ef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[675] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[676] = 80'h91b9a88b2186;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[676] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[677] = 80'hbaaaa92f9330;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[677] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[678] = 80'h899bc4d45fed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[678] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[679] = 80'h31aba86c07cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[679] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[680] = 80'hc4984e56b9a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[680] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[681] = 80'h1b2cb5378bd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[681] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[682] = 80'hff120ca68f9a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[682] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[683] = 80'ha835dfd4a64e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[683] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[684] = 80'hcc35683c57dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[684] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[685] = 80'ha5c1099a0ccc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[685] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[686] = 80'hefd95c4e5fe9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[686] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[687] = 80'h7c76d25796aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[687] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[688] = 80'h7b60730923d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[688] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[689] = 80'h7373b8b8f3c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[689] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[690] = 80'h37e56c799b77;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[690] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[691] = 80'h64aeec7ab84c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[691] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[692] = 80'hdc1814387312;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[692] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[693] = 80'hdd2835b8c4f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[693] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[694] = 80'h5af2eb552cca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[694] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[695] = 80'h446b9299fa74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[695] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[696] = 80'h86928cf64fc6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[696] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[697] = 80'hc4fdc019c61f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[697] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[698] = 80'h882f97bb161f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[698] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[699] = 80'h4ed606f4518d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[699] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem[700] = 80'hbd46a3aa3c15;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[0].u_tcam.mem_mask[700] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[1] = 80'h93d46a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[1] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[2] = 80'hd2356f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[2] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[3] = 80'h676259;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[3] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[4] = 80'h46079b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[4] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[5] = 80'h8c8892;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[5] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[6] = 80'h17cf44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[6] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[7] = 80'hbc724b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[7] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[8] = 80'he97981;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[8] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[9] = 80'h77a9de;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[9] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[10] = 80'h2b7a6c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[10] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[11] = 80'h504864;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[11] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[12] = 80'h8c6bb5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[12] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[13] = 80'h7afada;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[13] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[14] = 80'hcc3650;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[14] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[15] = 80'hdde1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[15] = 80'hffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[16] = 80'h41bae2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[16] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[17] = 80'h4b4f80;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[17] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[18] = 80'hccad23;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[18] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[19] = 80'h987d18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[19] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[20] = 80'h354214;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[20] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[21] = 80'h1b5bf0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[21] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[22] = 80'hcfcfe0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[22] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[23] = 80'h5dfdd7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[23] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[24] = 80'hf65193;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[24] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[25] = 80'h699932;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[25] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[26] = 80'h3c1356;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[26] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[27] = 80'hda35e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[27] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[28] = 80'hab08c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[28] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[29] = 80'h55162c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[29] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[30] = 80'h48ac99;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[30] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[31] = 80'hcf2b64;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[31] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[32] = 80'he09d8f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[32] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[33] = 80'h1d11e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[33] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[34] = 80'hdc6d6f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[34] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[35] = 80'h51d87e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[35] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[36] = 80'ha23c19;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[36] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[37] = 80'ha8d569;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[37] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[38] = 80'h9d9ed7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[38] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[39] = 80'h40e4d5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[39] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[40] = 80'h6b550f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[40] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[41] = 80'hb29e2e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[41] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[42] = 80'h2e7cf1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[42] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[43] = 80'h9200e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[43] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[44] = 80'hd9b933;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[44] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[45] = 80'hed726f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[45] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[46] = 80'h5a968d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[46] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[47] = 80'haa89df;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[47] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[48] = 80'hc1a0ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[48] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[49] = 80'h281727;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[49] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[50] = 80'hfe964b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[50] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[51] = 80'h649d6a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[51] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[52] = 80'hb66d0f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[52] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[53] = 80'ha77176;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[53] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[54] = 80'hab9e57;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[54] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[55] = 80'he15190;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[55] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[56] = 80'h935b3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[56] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[57] = 80'h7d3e7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[57] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[58] = 80'hd866b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[58] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[59] = 80'h4d2d96;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[59] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[60] = 80'h932137;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[60] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[61] = 80'hd76cda;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[61] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[62] = 80'hcfb810;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[62] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[63] = 80'h1f5e6f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[63] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[64] = 80'h866e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[64] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[65] = 80'h552409;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[65] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[66] = 80'h6819a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[66] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[67] = 80'hdabaa8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[67] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[68] = 80'h2fc8a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[68] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[69] = 80'h5014e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[69] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[70] = 80'hcc782f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[70] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[71] = 80'h6dae2a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[71] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[72] = 80'h39b496;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[72] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[73] = 80'h1cae91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[73] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[74] = 80'hcaff50;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[74] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[75] = 80'h33bd4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[75] = 80'h3ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[76] = 80'h4cb006;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[76] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[77] = 80'ha72599;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[77] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[78] = 80'h19efb1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[78] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[79] = 80'hbc0688;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[79] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[80] = 80'h37cb96;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[80] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[81] = 80'h65d77e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[81] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[82] = 80'ha4e182;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[82] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[83] = 80'hf9664b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[83] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[84] = 80'hd9d504;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[84] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[85] = 80'hac6429;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[85] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[86] = 80'h587b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[86] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[87] = 80'h70b9ff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[87] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[88] = 80'h7817b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[88] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[89] = 80'h5309c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[89] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[90] = 80'h263667;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[90] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[91] = 80'hbaef4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[91] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[92] = 80'h9fe398;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[92] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[93] = 80'hf404b2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[93] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[94] = 80'he66811;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[94] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[95] = 80'h6c4854;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[95] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[96] = 80'he41fbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[96] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[97] = 80'hae926c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[97] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[98] = 80'h8b4995;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[98] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[99] = 80'had9ee1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[99] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[100] = 80'he9cab6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[100] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[101] = 80'h190690;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[101] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[102] = 80'h644cd1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[102] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[103] = 80'h193143;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[103] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[104] = 80'hb38da9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[104] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[105] = 80'had42fb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[105] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[106] = 80'hf0c8e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[106] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[107] = 80'hc63e22;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[107] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[108] = 80'hceae4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[108] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[109] = 80'h81fce1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[109] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[110] = 80'h6c8b8a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[110] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[111] = 80'hc9c607;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[111] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[112] = 80'h84f36d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[112] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[113] = 80'h476c8a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[113] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[114] = 80'hd0a28d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[114] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[115] = 80'ha88374;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[115] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[116] = 80'hec0149;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[116] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[117] = 80'hd54c20;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[117] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[118] = 80'h990140;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[118] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[119] = 80'hd8c32b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[119] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[120] = 80'h9db7f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[120] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[121] = 80'h4fa872;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[121] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[122] = 80'hfa834c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[122] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[123] = 80'h640129;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[123] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[124] = 80'h472ab0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[124] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[125] = 80'hde8fce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[125] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[126] = 80'he5dd77;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[126] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[127] = 80'he2e528;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[127] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[128] = 80'hc4a88f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[128] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[129] = 80'h36d132;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[129] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[130] = 80'h103330;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[130] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[131] = 80'h210b4b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[131] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[132] = 80'h23a29c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[132] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[133] = 80'h18d134;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[133] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[134] = 80'h902d86;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[134] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[135] = 80'h599e1e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[135] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[136] = 80'h8b80f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[136] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[137] = 80'hfdd6d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[137] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[138] = 80'ha822ed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[138] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[139] = 80'h325c6b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[139] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[140] = 80'hf3a0f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[140] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[141] = 80'h40625f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[141] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[142] = 80'h62576;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[142] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[143] = 80'h247741;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[143] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[144] = 80'he66076;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[144] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[145] = 80'ha1bfdb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[145] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[146] = 80'h733a59;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[146] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[147] = 80'hd5364d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[147] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[148] = 80'hbf32c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[148] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[149] = 80'hdc5dbf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[149] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[150] = 80'h9a93fb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[150] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[151] = 80'hcf1ba8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[151] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[152] = 80'h2a29f0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[152] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[153] = 80'hdbde8b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[153] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[154] = 80'h9fe4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[154] = 80'hffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[155] = 80'h180c0a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[155] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[156] = 80'h88f835;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[156] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[157] = 80'h17109f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[157] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[158] = 80'h889713;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[158] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[159] = 80'h41b6b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[159] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[160] = 80'h864de9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[160] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[161] = 80'h7abce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[161] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[162] = 80'he12c35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[162] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[163] = 80'h301447;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[163] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[164] = 80'h76b32;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[164] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[165] = 80'h4b21b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[165] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[166] = 80'ha87adb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[166] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[167] = 80'h8e26bd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[167] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[168] = 80'he69464;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[168] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[169] = 80'hf1ae69;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[169] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[170] = 80'h3aec7a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[170] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[171] = 80'hee62e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[171] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[172] = 80'he8bc68;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[172] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[173] = 80'h5b86a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[173] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[174] = 80'h7871a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[174] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[175] = 80'h55f1d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[175] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[176] = 80'h96e694;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[176] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[177] = 80'h1fe63b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[177] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[178] = 80'h806547;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[178] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[179] = 80'h25c72f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[179] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[180] = 80'ha62af6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[180] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[181] = 80'h9d5417;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[181] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[182] = 80'h2c51af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[182] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[183] = 80'h2f7ca4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[183] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[184] = 80'hc3d2cf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[184] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[185] = 80'h2f8d88;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[185] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[186] = 80'h128302;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[186] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[187] = 80'h3cc6e7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[187] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[188] = 80'hbebdfb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[188] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[189] = 80'haaacbb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[189] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[190] = 80'h35afca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[190] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[191] = 80'h3f635d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[191] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[192] = 80'h9dc27f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[192] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[193] = 80'hf64438;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[193] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[194] = 80'h1cde19;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[194] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[195] = 80'had0b70;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[195] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[196] = 80'hb2a22c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[196] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[197] = 80'hc40815;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[197] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[198] = 80'ha08a15;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[198] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[199] = 80'h294352;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[199] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[200] = 80'h9f922;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[200] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[201] = 80'hc44933;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[201] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[202] = 80'hcba9fb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[202] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[203] = 80'hcee397;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[203] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[204] = 80'h5ab855;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[204] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[205] = 80'hc37cff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[205] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[206] = 80'hf1815;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[206] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[207] = 80'h1fecf8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[207] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[208] = 80'h2f0cd3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[208] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[209] = 80'hcdfdc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[209] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[210] = 80'heada3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[210] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[211] = 80'hc5239f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[211] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[212] = 80'h2e0306;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[212] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[213] = 80'h9b50e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[213] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[214] = 80'h244d2d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[214] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[215] = 80'hd04cf1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[215] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[216] = 80'h12056a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[216] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[217] = 80'h17ca62;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[217] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[218] = 80'h3f7a75;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[218] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[219] = 80'h7a839f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[219] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[220] = 80'h488d5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[220] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[221] = 80'h34ae81;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[221] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[222] = 80'h1ee202;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[222] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[223] = 80'h183ea5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[223] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[224] = 80'hc5cf43;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[224] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[225] = 80'he2bc13;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[225] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[226] = 80'h1fd051;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[226] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[227] = 80'h1d970f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[227] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[228] = 80'hc403c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[228] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[229] = 80'h88f8af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[229] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[230] = 80'h522f39;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[230] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[231] = 80'hf385d1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[231] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[232] = 80'h9777c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[232] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[233] = 80'hffee98;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[233] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[234] = 80'h8f8852;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[234] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[235] = 80'h22a823;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[235] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[236] = 80'haabbdd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[236] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[237] = 80'hc4d792;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[237] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[238] = 80'h1af82d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[238] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[239] = 80'h12e62a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[239] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[240] = 80'h84feb8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[240] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[241] = 80'he90935;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[241] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[242] = 80'hdaeacf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[242] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[243] = 80'hf7fb36;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[243] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[244] = 80'hb754c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[244] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[245] = 80'h72a0d2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[245] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[246] = 80'h14c7a8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[246] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[247] = 80'h2e7ccb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[247] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[248] = 80'h172d6b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[248] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[249] = 80'h5cbd69;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[249] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[250] = 80'h838848;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[250] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[251] = 80'he57f48;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[251] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[252] = 80'h879954;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[252] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[253] = 80'h3f3b48;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[253] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[254] = 80'haa15a1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[254] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[255] = 80'h72e889;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[255] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[256] = 80'h1b542;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[256] = 80'h1ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[257] = 80'h296632;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[257] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[258] = 80'h38ad9e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[258] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[259] = 80'hdd5b20;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[259] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[260] = 80'h7e3d3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[260] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[261] = 80'hde577e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[261] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[262] = 80'h5f90c0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[262] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[263] = 80'hd30cb2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[263] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[264] = 80'h8ebe76;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[264] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[265] = 80'h2d1e33;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[265] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[266] = 80'h78e2fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[266] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[267] = 80'h8595a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[267] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[268] = 80'h4d7b60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[268] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[269] = 80'ha5d4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[269] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[270] = 80'hb6a7b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[270] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[271] = 80'hb9d0d8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[271] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[272] = 80'h7c54d0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[272] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[273] = 80'hfab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[273] = 80'hfff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[274] = 80'h526452;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[274] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[275] = 80'heea715;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[275] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[276] = 80'hb958bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[276] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[277] = 80'ha9b50c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[277] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[278] = 80'hfcbf5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[278] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[279] = 80'hd7128e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[279] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[280] = 80'h287b14;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[280] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[281] = 80'h99d893;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[281] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[282] = 80'hce1be7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[282] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[283] = 80'h275c14;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[283] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[284] = 80'hb2ecf6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[284] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[285] = 80'h32209f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[285] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[286] = 80'h8890e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[286] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[287] = 80'h5df3a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[287] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[288] = 80'h681f7e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[288] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[289] = 80'h52ac42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[289] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[290] = 80'h62b76d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[290] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[291] = 80'h2a3054;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[291] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[292] = 80'ha6aacb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[292] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[293] = 80'hfad7b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[293] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[294] = 80'he45af7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[294] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[295] = 80'h1b8312;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[295] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[296] = 80'h4d7686;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[296] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[297] = 80'h9e9f11;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[297] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[298] = 80'h3752b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[298] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[299] = 80'h9fff19;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[299] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[300] = 80'h3deeb0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[300] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[301] = 80'h4d0cc0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[301] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[302] = 80'had4e0b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[302] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[303] = 80'hd93c76;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[303] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[304] = 80'ha363f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[304] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[305] = 80'hfe7a4a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[305] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[306] = 80'h6750fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[306] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[307] = 80'hfa4199;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[307] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[308] = 80'hd91f85;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[308] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[309] = 80'h6021c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[309] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[310] = 80'hb7fc65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[310] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[311] = 80'hd6e41;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[311] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[312] = 80'h1fc6a1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[312] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[313] = 80'hd152b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[313] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[314] = 80'h2f8780;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[314] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[315] = 80'ha9948;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[315] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[316] = 80'h249ab8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[316] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[317] = 80'h472875;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[317] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[318] = 80'h6d2196;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[318] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[319] = 80'h10373f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[319] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[320] = 80'hc0f50e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[320] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[321] = 80'hdd84a8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[321] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[322] = 80'h324444;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[322] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[323] = 80'hb11fe3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[323] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[324] = 80'hd3c003;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[324] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[325] = 80'h22c068;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[325] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[326] = 80'h200557;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[326] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[327] = 80'hd760d5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[327] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[328] = 80'h404d84;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[328] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[329] = 80'h38a6a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[329] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[330] = 80'h3a4640;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[330] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[331] = 80'h4a10b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[331] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[332] = 80'hb30115;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[332] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[333] = 80'h8aeaa5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[333] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[334] = 80'hf1cc59;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[334] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[335] = 80'h7f6f35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[335] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[336] = 80'h465838;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[336] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[337] = 80'hc08db5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[337] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[338] = 80'hfd7be1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[338] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[339] = 80'ha0f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[339] = 80'hffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[340] = 80'hb91869;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[340] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[341] = 80'hc0ad63;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[341] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[342] = 80'hb08e22;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[342] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[343] = 80'hf68553;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[343] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[344] = 80'h64927f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[344] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[345] = 80'h83a02e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[345] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[346] = 80'hbe5a96;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[346] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[347] = 80'h6e40d1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[347] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[348] = 80'hf76daa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[348] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[349] = 80'h260806;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[349] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[350] = 80'haaf348;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[350] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[351] = 80'hbe1a7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[351] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[352] = 80'ha59283;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[352] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[353] = 80'h9fd1ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[353] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[354] = 80'h8acbff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[354] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[355] = 80'h4deca7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[355] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[356] = 80'h28e13a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[356] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[357] = 80'ha299ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[357] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[358] = 80'h99a477;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[358] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[359] = 80'h44a766;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[359] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[360] = 80'hd3a394;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[360] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[361] = 80'hecc3e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[361] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[362] = 80'hebab0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[362] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[363] = 80'h7f07a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[363] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[364] = 80'h1940da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[364] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[365] = 80'hdd77fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[365] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[366] = 80'h27a422;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[366] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[367] = 80'he19559;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[367] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[368] = 80'h8d63;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[368] = 80'hffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[369] = 80'h1193c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[369] = 80'h1ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[370] = 80'h46a7c0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[370] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[371] = 80'hc71745;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[371] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[372] = 80'hee0321;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[372] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[373] = 80'h21c943;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[373] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[374] = 80'h5334c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[374] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[375] = 80'hcbd414;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[375] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[376] = 80'hab0538;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[376] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[377] = 80'hf176c0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[377] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[378] = 80'h8512ed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[378] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[379] = 80'ha0128d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[379] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[380] = 80'hdb3124;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[380] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[381] = 80'h3d7888;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[381] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[382] = 80'h6f91b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[382] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[383] = 80'hb21e43;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[383] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[384] = 80'h8de00c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[384] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[385] = 80'had6a91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[385] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[386] = 80'h9982b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[386] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[387] = 80'hf936b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[387] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[388] = 80'hfb8434;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[388] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[389] = 80'h61ac31;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[389] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[390] = 80'hd66;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[390] = 80'hfff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[391] = 80'hcb4d6b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[391] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[392] = 80'h952555;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[392] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[393] = 80'hd662de;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[393] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[394] = 80'haa0ea6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[394] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[395] = 80'hba2e0f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[395] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[396] = 80'hf7491c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[396] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[397] = 80'h8d68ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[397] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[398] = 80'ha366a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[398] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[399] = 80'h7672fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[399] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[400] = 80'h4e0e5b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[400] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[401] = 80'hf69f93;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[401] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[402] = 80'hdc64a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[402] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[403] = 80'h3e36d7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[403] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[404] = 80'h20cd14;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[404] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[405] = 80'hfd80ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[405] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[406] = 80'h14a853;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[406] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[407] = 80'hd34e71;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[407] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[408] = 80'h4da43e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[408] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[409] = 80'h2dcdd0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[409] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[410] = 80'hff51e4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[410] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[411] = 80'h5e4c3b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[411] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[412] = 80'h919a50;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[412] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[413] = 80'h5c6f6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[413] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[414] = 80'h4880e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[414] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[415] = 80'hb52f6e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[415] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[416] = 80'h6330f5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[416] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[417] = 80'h87589c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[417] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[418] = 80'hae87c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[418] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[419] = 80'h88b591;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[419] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[420] = 80'ha9681c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[420] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[421] = 80'h5bfe8c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[421] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[422] = 80'hfeeabb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[422] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[423] = 80'h5bfef3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[423] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[424] = 80'hc439f5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[424] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[425] = 80'hcbb611;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[425] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[426] = 80'h6bf841;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[426] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[427] = 80'h14eb96;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[427] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[428] = 80'hcb6ce3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[428] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[429] = 80'hbe0907;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[429] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[430] = 80'hf515b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[430] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[431] = 80'hd4b21b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[431] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[432] = 80'haed1b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[432] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[433] = 80'h187e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[433] = 80'h1ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[434] = 80'h3bf896;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[434] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[435] = 80'hd53055;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[435] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[436] = 80'hd85a46;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[436] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[437] = 80'hb70da5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[437] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[438] = 80'hf14efb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[438] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[439] = 80'hceed54;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[439] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[440] = 80'h1c63cc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[440] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[441] = 80'h2e657b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[441] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[442] = 80'h1b7bb1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[442] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[443] = 80'ha490bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[443] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[444] = 80'h77f7c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[444] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[445] = 80'hce3879;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[445] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[446] = 80'h3d62f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[446] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[447] = 80'hd3c317;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[447] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[448] = 80'hcd4052;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[448] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[449] = 80'h366029;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[449] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[450] = 80'h249c31;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[450] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[451] = 80'hf85353;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[451] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[452] = 80'hba861d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[452] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[453] = 80'h7b4f14;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[453] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[454] = 80'he9a8b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[454] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[455] = 80'h48daff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[455] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[456] = 80'h9eeb3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[456] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[457] = 80'h1ea67;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[457] = 80'h1ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[458] = 80'hb2c532;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[458] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[459] = 80'h8cdabd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[459] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[460] = 80'he33611;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[460] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[461] = 80'h888646;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[461] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[462] = 80'h7532ec;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[462] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[463] = 80'hef77eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[463] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[464] = 80'h836a74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[464] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[465] = 80'h60abde;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[465] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[466] = 80'h1fb207;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[466] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[467] = 80'h1fd4bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[467] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[468] = 80'he37673;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[468] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[469] = 80'he78f3e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[469] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[470] = 80'hf089bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[470] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[471] = 80'h989a46;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[471] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[472] = 80'h4872d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[472] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[473] = 80'h7d4a59;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[473] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[474] = 80'h79148c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[474] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[475] = 80'hca4d53;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[475] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[476] = 80'h318859;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[476] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[477] = 80'hd19af7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[477] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[478] = 80'h270545;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[478] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[479] = 80'h94a8f5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[479] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[480] = 80'hfd4a65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[480] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[481] = 80'h14a4ed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[481] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[482] = 80'hb279ba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[482] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[483] = 80'h63905b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[483] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[484] = 80'h528285;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[484] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[485] = 80'hbd6eb1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[485] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[486] = 80'h136e6c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[486] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[487] = 80'h9b3456;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[487] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[488] = 80'h254c0a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[488] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[489] = 80'hec438c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[489] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[490] = 80'h84699d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[490] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[491] = 80'hd0224;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[491] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[492] = 80'hc49916;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[492] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[493] = 80'hff4173;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[493] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[494] = 80'h81bccf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[494] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[495] = 80'h6fed17;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[495] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[496] = 80'h2329d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[496] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[497] = 80'he35295;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[497] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[498] = 80'h97a6ce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[498] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[499] = 80'h7355fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[499] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[500] = 80'hb5e794;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[500] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[501] = 80'h3295ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[501] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[502] = 80'heca5ce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[502] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[503] = 80'h87bf14;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[503] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[504] = 80'ha166f5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[504] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[505] = 80'hc0b98a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[505] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[506] = 80'h452cdc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[506] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[507] = 80'h78e1e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[507] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[508] = 80'h92eb8c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[508] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[509] = 80'h129629;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[509] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[510] = 80'hbc837b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[510] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[511] = 80'h9cda8f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[511] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[512] = 80'h3e36f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[512] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[513] = 80'h8a27cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[513] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[514] = 80'h462c62;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[514] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[515] = 80'hdfcade;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[515] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[516] = 80'h8989c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[516] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[517] = 80'h6c0294;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[517] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[518] = 80'hbcd2eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[518] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[519] = 80'h3bff68;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[519] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[520] = 80'h6b9b27;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[520] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[521] = 80'h22b3ea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[521] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[522] = 80'h41688a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[522] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[523] = 80'he21345;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[523] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[524] = 80'h73d32b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[524] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[525] = 80'ha2a953;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[525] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[526] = 80'h4e430c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[526] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[527] = 80'h64d84c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[527] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[528] = 80'h2f0b4c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[528] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[529] = 80'h3b69f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[529] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[530] = 80'hac0c0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[530] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[531] = 80'h2cb8c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[531] = 80'h3ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[532] = 80'hc8973d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[532] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[533] = 80'h63403b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[533] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[534] = 80'h3b10ba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[534] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[535] = 80'h2ce7ba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[535] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[536] = 80'hea87;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[536] = 80'hffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[537] = 80'h50badf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[537] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[538] = 80'h5b2fbb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[538] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[539] = 80'hac32d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[539] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[540] = 80'h175207;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[540] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[541] = 80'hce27f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[541] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[542] = 80'h75d740;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[542] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[543] = 80'h76d79a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[543] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[544] = 80'h7390f8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[544] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[545] = 80'hb963bf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[545] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[546] = 80'h26405;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[546] = 80'h3ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[547] = 80'ha04b21;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[547] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[548] = 80'ha30541;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[548] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[549] = 80'h8927b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[549] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[550] = 80'h9cc1c0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[550] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[551] = 80'h3ba3f5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[551] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[552] = 80'h352e1d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[552] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[553] = 80'hc2fbc1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[553] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[554] = 80'h4cbb09;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[554] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[555] = 80'hffbbbf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[555] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[556] = 80'hb682c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[556] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[557] = 80'h52c4da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[557] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[558] = 80'h312a41;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[558] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[559] = 80'h8b4d5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[559] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[560] = 80'hf3a2ad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[560] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[561] = 80'h6e7c4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[561] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[562] = 80'hded8dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[562] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[563] = 80'h1dc81;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[563] = 80'h1ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[564] = 80'hfbaf9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[564] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[565] = 80'h61584b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[565] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[566] = 80'h7649b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[566] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[567] = 80'h5f5cd1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[567] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[568] = 80'hf10131;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[568] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[569] = 80'h72671c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[569] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[570] = 80'hd3785d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[570] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[571] = 80'ha29593;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[571] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[572] = 80'h954c60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[572] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[573] = 80'hc17e8e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[573] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[574] = 80'h9a7ba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[574] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[575] = 80'h7072f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[575] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[576] = 80'h78fcbf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[576] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[577] = 80'h43c1b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[577] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[578] = 80'hb08007;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[578] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[579] = 80'h150566;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[579] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[580] = 80'ha9a978;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[580] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[581] = 80'hc86b86;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[581] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[582] = 80'hf6a9b4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[582] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[583] = 80'hbd5e1d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[583] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[584] = 80'h6bdf3d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[584] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[585] = 80'h8848ec;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[585] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[586] = 80'h2de4cb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[586] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[587] = 80'h729081;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[587] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[588] = 80'h6a8d3d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[588] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[589] = 80'hb986e7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[589] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[590] = 80'h53a9dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[590] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[591] = 80'h495aab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[591] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[592] = 80'h2243c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[592] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[593] = 80'h932bc5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[593] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[594] = 80'hc7e5a1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[594] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[595] = 80'h519f51;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[595] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[596] = 80'h31d9d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[596] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[597] = 80'h6c648c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[597] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[598] = 80'hca4098;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[598] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[599] = 80'he6aa63;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[599] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[600] = 80'h9898d6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[600] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[601] = 80'h2e0ee6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[601] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[602] = 80'h7de959;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[602] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[603] = 80'h22ed5e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[603] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[604] = 80'hef9cd4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[604] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[605] = 80'h9e573b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[605] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[606] = 80'ha4a6bf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[606] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[607] = 80'h96fae7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[607] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[608] = 80'hcdbaec;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[608] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[609] = 80'hf9a463;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[609] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[610] = 80'h4e36e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[610] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[611] = 80'hf0a7a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[611] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[612] = 80'h1ae7e7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[612] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[613] = 80'hfacdcc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[613] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[614] = 80'h57f90;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[614] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[615] = 80'hb782da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[615] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[616] = 80'h68b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[616] = 80'h7fff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[617] = 80'h3a8542;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[617] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[618] = 80'h662a36;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[618] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[619] = 80'hc447e7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[619] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[620] = 80'h428275;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[620] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[621] = 80'h207e9f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[621] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[622] = 80'hb5de9b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[622] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[623] = 80'hbdfb18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[623] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[624] = 80'h3a7a85;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[624] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[625] = 80'h6b085d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[625] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[626] = 80'he56816;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[626] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[627] = 80'h18d22b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[627] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[628] = 80'hfd73c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[628] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[629] = 80'hf65166;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[629] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[630] = 80'haea4f6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[630] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[631] = 80'h378ad7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[631] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[632] = 80'h7215cb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[632] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[633] = 80'h4370d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[633] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[634] = 80'he0bb48;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[634] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[635] = 80'hdd2dbc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[635] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[636] = 80'hd10c0d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[636] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[637] = 80'h45ca7b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[637] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[638] = 80'h50ec64;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[638] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[639] = 80'h906144;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[639] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[640] = 80'h112dc1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[640] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[641] = 80'h5b36ae;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[641] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[642] = 80'h6a5c37;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[642] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[643] = 80'h24a942;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[643] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[644] = 80'h48e2b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[644] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[645] = 80'h77fa27;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[645] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[646] = 80'h78b151;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[646] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[647] = 80'ha47604;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[647] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[648] = 80'h594a3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[648] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[649] = 80'haf2e91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[649] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[650] = 80'h54f406;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[650] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[651] = 80'hdbd353;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[651] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[652] = 80'ha961f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[652] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[653] = 80'h655384;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[653] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[654] = 80'h1b8b2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[654] = 80'h1ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[655] = 80'hb646a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[655] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[656] = 80'hc35541;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[656] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[657] = 80'haa459d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[657] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[658] = 80'h759b4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[658] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[659] = 80'h10b764;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[659] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[660] = 80'h7f2ca2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[660] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[661] = 80'h9605;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[661] = 80'hffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[662] = 80'h880ee7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[662] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[663] = 80'heced99;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[663] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[664] = 80'h8a05ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[664] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[665] = 80'h66baf9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[665] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[666] = 80'h96805d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[666] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[667] = 80'he3de2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[667] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[668] = 80'h15e3df;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[668] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[669] = 80'ha47712;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[669] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[670] = 80'h1932f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[670] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[671] = 80'h15d54c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[671] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[672] = 80'h8e6097;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[672] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[673] = 80'h26723;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[673] = 80'h3ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[674] = 80'h2d4201;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[674] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[675] = 80'h64a019;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[675] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[676] = 80'h52068;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[676] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[677] = 80'h4fc87f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[677] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[678] = 80'h354c4a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[678] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[679] = 80'hc084df;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[679] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[680] = 80'he3af6c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[680] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[681] = 80'h9b4c6a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[681] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[682] = 80'h4fe061;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[682] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[683] = 80'h668b54;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[683] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[684] = 80'hb7d2fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[684] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[685] = 80'h7b394b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[685] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[686] = 80'ha0d693;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[686] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[687] = 80'hecb9e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[687] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[688] = 80'hfa6dcb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[688] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[689] = 80'h549727;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[689] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[690] = 80'h563be7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[690] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[691] = 80'hefc0f2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[691] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[692] = 80'hc5e4f2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[692] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[693] = 80'h97e2e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[693] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[694] = 80'hd71d42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[694] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[695] = 80'h2cc08f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[695] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[696] = 80'h6e18f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[696] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[697] = 80'hfdf59;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[697] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[698] = 80'h8f22b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[698] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[699] = 80'hf70e50;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[699] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem[700] = 80'h65c364;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[3].u_tcam.mem_mask[700] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[1] = 80'h7f1ea9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[1] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[2] = 80'h18d7d4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[2] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[3] = 80'h879503;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[3] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[4] = 80'h795e9d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[4] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[5] = 80'hd8811f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[5] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[6] = 80'hf72c4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[6] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[7] = 80'h45bc37;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[7] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[8] = 80'ha9ca1e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[8] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[9] = 80'h95fadc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[9] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[10] = 80'hfd7856;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[10] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[11] = 80'h3ac1d0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[11] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[12] = 80'hc47e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[12] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[13] = 80'hfb27f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[13] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[14] = 80'h18fca4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[14] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[15] = 80'h2e4356;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[15] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[16] = 80'h56a40c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[16] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[17] = 80'h18540e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[17] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[18] = 80'hea2b44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[18] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[19] = 80'h84c769;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[19] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[20] = 80'h9ae0b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[20] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[21] = 80'ha15356;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[21] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[22] = 80'h5a0605;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[22] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[23] = 80'h6fe0cb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[23] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[24] = 80'he646d6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[24] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[25] = 80'ha2d6b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[25] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[26] = 80'hf04d5b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[26] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[27] = 80'h4c578c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[27] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[28] = 80'h888d1f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[28] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[29] = 80'h2ca3fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[29] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[30] = 80'h63455b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[30] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[31] = 80'h2768c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[31] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[32] = 80'h7cb8cb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[32] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[33] = 80'h62f735;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[33] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[34] = 80'h2fa2ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[34] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[35] = 80'h6b0b30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[35] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[36] = 80'hdc4120;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[36] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[37] = 80'hd471aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[37] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[38] = 80'h40a7fc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[38] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[39] = 80'hac33c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[39] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[40] = 80'h109775;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[40] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[41] = 80'hc3ff40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[41] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[42] = 80'h283e24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[42] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[43] = 80'hd2bca2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[43] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[44] = 80'h5178a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[44] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[45] = 80'h9ab1a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[45] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[46] = 80'hdd0418;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[46] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[47] = 80'h4341e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[47] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[48] = 80'hbeafd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[48] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[49] = 80'h653c68;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[49] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[50] = 80'hc2f7fb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[50] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[51] = 80'h2ec425;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[51] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[52] = 80'h39f1b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[52] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[53] = 80'h65b81f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[53] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[54] = 80'he84bff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[54] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[55] = 80'h6f12c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[55] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[56] = 80'h638539;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[56] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[57] = 80'h74386b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[57] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[58] = 80'h6ec296;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[58] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[59] = 80'h9dc45a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[59] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[60] = 80'h7bdeb2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[60] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[61] = 80'h109400;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[61] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[62] = 80'h3ed34b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[62] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[63] = 80'h83a39a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[63] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[64] = 80'hb39350;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[64] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[65] = 80'h3fd68e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[65] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[66] = 80'h168dc8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[66] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[67] = 80'hc7d864;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[67] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[68] = 80'h6ac4b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[68] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[69] = 80'h29c5fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[69] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[70] = 80'h7775e4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[70] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[71] = 80'h354a38;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[71] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[72] = 80'h482f82;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[72] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[73] = 80'h8f4dc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[73] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[74] = 80'h2f794e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[74] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[75] = 80'hc688bd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[75] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[76] = 80'h8c6bf8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[76] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[77] = 80'h4a580d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[77] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[78] = 80'he51d07;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[78] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[79] = 80'h6576cb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[79] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[80] = 80'h672b33;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[80] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[81] = 80'h765369;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[81] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[82] = 80'h65548;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[82] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[83] = 80'hfa8b7f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[83] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[84] = 80'h9e0149;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[84] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[85] = 80'h3700bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[85] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[86] = 80'ha26d54;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[86] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[87] = 80'h485e50;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[87] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[88] = 80'h4e377c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[88] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[89] = 80'h290bd8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[89] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[90] = 80'h79eac3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[90] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[91] = 80'haeb963;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[91] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[92] = 80'he60f6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[92] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[93] = 80'hebc64c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[93] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[94] = 80'hfd79da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[94] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[95] = 80'h5f903f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[95] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[96] = 80'h8c6098;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[96] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[97] = 80'h52bbf8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[97] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[98] = 80'h67064a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[98] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[99] = 80'heda0ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[99] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[100] = 80'h9fe0b2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[100] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[101] = 80'h2b0b9e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[101] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[102] = 80'h8ed315;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[102] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[103] = 80'h3fa5eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[103] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[104] = 80'hd5a9ea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[104] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[105] = 80'h3b5063;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[105] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[106] = 80'h3de498;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[106] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[107] = 80'h34d05b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[107] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[108] = 80'h9906b4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[108] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[109] = 80'h8e8559;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[109] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[110] = 80'he3f52;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[110] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[111] = 80'h4b4571;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[111] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[112] = 80'h1da95e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[112] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[113] = 80'hf8a77d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[113] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[114] = 80'h773e7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[114] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[115] = 80'hcc18d8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[115] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[116] = 80'h523f2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[116] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[117] = 80'hd32eb1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[117] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[118] = 80'hb10a04;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[118] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[119] = 80'h9e289a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[119] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[120] = 80'h3f745c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[120] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[121] = 80'hb4d716;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[121] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[122] = 80'h353aba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[122] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[123] = 80'h138266;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[123] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[124] = 80'h98c3a8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[124] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[125] = 80'ha72bb0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[125] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[126] = 80'hf0a808;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[126] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[127] = 80'h2ecc7c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[127] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[128] = 80'h70432e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[128] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[129] = 80'h9e5629;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[129] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[130] = 80'hb9028f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[130] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[131] = 80'h7d192f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[131] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[132] = 80'h9f9291;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[132] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[133] = 80'hee6a20;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[133] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[134] = 80'h53672d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[134] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[135] = 80'hdd027c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[135] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[136] = 80'hdc08c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[136] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[137] = 80'h58402c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[137] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[138] = 80'hc81a4a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[138] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[139] = 80'hedd5d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[139] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[140] = 80'h4b52;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[140] = 80'h7fff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[141] = 80'he03ed4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[141] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[142] = 80'h7e9436;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[142] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[143] = 80'h784bef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[143] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[144] = 80'h42f39d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[144] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[145] = 80'hbe6a7e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[145] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[146] = 80'h826f57;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[146] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[147] = 80'h29e2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[147] = 80'h3ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[148] = 80'h29c960;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[148] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[149] = 80'h19c756;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[149] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[150] = 80'h1fbdf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[150] = 80'h1ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[151] = 80'h798a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[151] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[152] = 80'h376c99;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[152] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[153] = 80'h2e7c93;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[153] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[154] = 80'h6e0c48;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[154] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[155] = 80'h7848e4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[155] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[156] = 80'heab49b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[156] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[157] = 80'h3c4183;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[157] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[158] = 80'h206e77;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[158] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[159] = 80'h60af7b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[159] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[160] = 80'h532847;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[160] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[161] = 80'hbad608;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[161] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[162] = 80'h47a19a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[162] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[163] = 80'hf8c422;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[163] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[164] = 80'h9c50ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[164] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[165] = 80'h2c4a16;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[165] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[166] = 80'he2f212;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[166] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[167] = 80'h32b6e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[167] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[168] = 80'h501cd9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[168] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[169] = 80'h59d817;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[169] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[170] = 80'h79c4b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[170] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[171] = 80'hdbfb38;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[171] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[172] = 80'h3c8d91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[172] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[173] = 80'h700b97;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[173] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[174] = 80'h6a6798;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[174] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[175] = 80'hb16541;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[175] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[176] = 80'h148fdc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[176] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[177] = 80'hc77ae0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[177] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[178] = 80'h289a41;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[178] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[179] = 80'hcce9c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[179] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[180] = 80'h3293d0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[180] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[181] = 80'h85fe27;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[181] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[182] = 80'h7de321;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[182] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[183] = 80'h556878;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[183] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[184] = 80'ha2e200;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[184] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[185] = 80'hf7b199;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[185] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[186] = 80'h4e7d0f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[186] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[187] = 80'h2932d5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[187] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[188] = 80'hf10ee2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[188] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[189] = 80'hd3cb30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[189] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[190] = 80'hdc4082;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[190] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[191] = 80'h4680df;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[191] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[192] = 80'h3e3ace;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[192] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[193] = 80'h278237;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[193] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[194] = 80'hf58b4b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[194] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[195] = 80'h53a60b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[195] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[196] = 80'h29bce4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[196] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[197] = 80'hbf1a0a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[197] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[198] = 80'he19318;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[198] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[199] = 80'h44d266;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[199] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[200] = 80'ha6b455;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[200] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[201] = 80'ha1ed9d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[201] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[202] = 80'h4fc0f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[202] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[203] = 80'h83eaaf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[203] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[204] = 80'h1d8f2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[204] = 80'h1ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[205] = 80'hc8461;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[205] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[206] = 80'h5a9ad8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[206] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[207] = 80'h45adc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[207] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[208] = 80'h44e7f5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[208] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[209] = 80'h4a5dba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[209] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[210] = 80'h82d37a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[210] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[211] = 80'ha5936e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[211] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[212] = 80'h7b239;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[212] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[213] = 80'h12fd45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[213] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[214] = 80'h842ec1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[214] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[215] = 80'h5fee07;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[215] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[216] = 80'h386dc0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[216] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[217] = 80'h30a003;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[217] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[218] = 80'h69dabf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[218] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[219] = 80'hc8cd9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[219] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[220] = 80'h20926d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[220] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[221] = 80'hc358af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[221] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[222] = 80'h5bb9eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[222] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[223] = 80'hb1e73e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[223] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[224] = 80'h591f46;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[224] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[225] = 80'h7367d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[225] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[226] = 80'h638b62;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[226] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[227] = 80'h637b90;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[227] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[228] = 80'h8d74b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[228] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[229] = 80'h5c8f52;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[229] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[230] = 80'hd7ee49;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[230] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[231] = 80'hd72b91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[231] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[232] = 80'h816c24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[232] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[233] = 80'hde97a8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[233] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[234] = 80'h4ef26b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[234] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[235] = 80'hafbc7c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[235] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[236] = 80'h337d7d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[236] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[237] = 80'h781a2b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[237] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[238] = 80'hb4e99c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[238] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[239] = 80'ha1d931;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[239] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[240] = 80'h2e3027;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[240] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[241] = 80'hf983f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[241] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[242] = 80'h56ed80;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[242] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[243] = 80'h5200ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[243] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[244] = 80'h637797;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[244] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[245] = 80'hdd2137;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[245] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[246] = 80'hfd2416;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[246] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[247] = 80'hf3a4f0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[247] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[248] = 80'h44c886;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[248] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[249] = 80'hceb410;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[249] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[250] = 80'hf59b12;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[250] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[251] = 80'he49bd0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[251] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[252] = 80'h638997;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[252] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[253] = 80'h2f7580;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[253] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[254] = 80'h1c10a8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[254] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[255] = 80'h879f04;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[255] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[256] = 80'hbab2c4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[256] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[257] = 80'ha22715;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[257] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[258] = 80'hf23b5e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[258] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[259] = 80'hfdc001;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[259] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[260] = 80'h288bf0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[260] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[261] = 80'h662d40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[261] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[262] = 80'h72cef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[262] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[263] = 80'h87666;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[263] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[264] = 80'hf522c4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[264] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[265] = 80'hcf63c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[265] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[266] = 80'he18e89;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[266] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[267] = 80'ha2bc46;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[267] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[268] = 80'h41996f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[268] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[269] = 80'h5e2a51;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[269] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[270] = 80'h46b451;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[270] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[271] = 80'hee2aae;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[271] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[272] = 80'hb33948;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[272] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[273] = 80'h7587fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[273] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[274] = 80'h4584c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[274] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[275] = 80'h4532c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[275] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[276] = 80'h7754d8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[276] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[277] = 80'h2b77b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[277] = 80'h3ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[278] = 80'h8f7473;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[278] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[279] = 80'hff2471;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[279] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[280] = 80'h14b05f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[280] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[281] = 80'hdf9570;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[281] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[282] = 80'h153dbb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[282] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[283] = 80'hc5d62c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[283] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[284] = 80'h6bf1fb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[284] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[285] = 80'h25d7ea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[285] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[286] = 80'h7d1082;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[286] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[287] = 80'h5f39c9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[287] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[288] = 80'h9fe99;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[288] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[289] = 80'h7b04db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[289] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[290] = 80'h29dd6a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[290] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[291] = 80'h1fcd7e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[291] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[292] = 80'h5b635c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[292] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[293] = 80'h6eda0f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[293] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[294] = 80'hcef008;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[294] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[295] = 80'h32dc5e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[295] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[296] = 80'h50586f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[296] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[297] = 80'h6dc367;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[297] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[298] = 80'h9c1de1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[298] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[299] = 80'hfd77d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[299] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[300] = 80'hd3c5d4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[300] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[301] = 80'hfdb0d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[301] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[302] = 80'h25d51;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[302] = 80'h3ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[303] = 80'he88800;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[303] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[304] = 80'hc08b8e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[304] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[305] = 80'h3f0392;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[305] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[306] = 80'ha02fb5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[306] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[307] = 80'h21607f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[307] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[308] = 80'h8f612f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[308] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[309] = 80'h34a36e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[309] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[310] = 80'h899446;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[310] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[311] = 80'haeaee1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[311] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[312] = 80'hefa58;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[312] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[313] = 80'h7c121d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[313] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[314] = 80'h84c243;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[314] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[315] = 80'h6fa6f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[315] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[316] = 80'he50d93;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[316] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[317] = 80'h30a2f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[317] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[318] = 80'h28773f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[318] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[319] = 80'h266b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[319] = 80'h3ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[320] = 80'ha9817d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[320] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[321] = 80'h3920db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[321] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[322] = 80'h3bfaad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[322] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[323] = 80'hd9c7f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[323] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[324] = 80'h5c0486;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[324] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[325] = 80'hd00200;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[325] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[326] = 80'hd49869;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[326] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[327] = 80'h89ee4e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[327] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[328] = 80'hdf942f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[328] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[329] = 80'h84601d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[329] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[330] = 80'h1808be;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[330] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[331] = 80'hb502fb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[331] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[332] = 80'h9f2b20;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[332] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[333] = 80'hb2fa64;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[333] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[334] = 80'h80dd3b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[334] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[335] = 80'h38568a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[335] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[336] = 80'hea6666;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[336] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[337] = 80'hdfa001;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[337] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[338] = 80'h396ef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[338] = 80'h3ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[339] = 80'h61ba43;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[339] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[340] = 80'h80209;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[340] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[341] = 80'h5b8fa1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[341] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[342] = 80'h61c5cc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[342] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[343] = 80'hb26ef1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[343] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[344] = 80'h407501;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[344] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[345] = 80'h28ace5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[345] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[346] = 80'hc579b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[346] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[347] = 80'h9bfb01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[347] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[348] = 80'hf34eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[348] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[349] = 80'hab2f3d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[349] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[350] = 80'h186408;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[350] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[351] = 80'h22a3c9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[351] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[352] = 80'h9aa041;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[352] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[353] = 80'hb46f64;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[353] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[354] = 80'h48548b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[354] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[355] = 80'he7ee30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[355] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[356] = 80'hc7e65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[356] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[357] = 80'hc4e05f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[357] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[358] = 80'hcdeb94;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[358] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[359] = 80'hc6fbde;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[359] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[360] = 80'h4364d2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[360] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[361] = 80'h54c878;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[361] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[362] = 80'h244700;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[362] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[363] = 80'h3a7f6d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[363] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[364] = 80'he03a58;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[364] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[365] = 80'hb0efa4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[365] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[366] = 80'h1e6831;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[366] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[367] = 80'h323acf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[367] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[368] = 80'h1ab23b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[368] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[369] = 80'h153918;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[369] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[370] = 80'ha376d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[370] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[371] = 80'h66c250;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[371] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[372] = 80'hf46295;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[372] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[373] = 80'h909a33;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[373] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[374] = 80'hb903f6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[374] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[375] = 80'h876713;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[375] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[376] = 80'hf203b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[376] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[377] = 80'h7035e4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[377] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[378] = 80'he24033;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[378] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[379] = 80'he8a4a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[379] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[380] = 80'hece548;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[380] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[381] = 80'h586dfc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[381] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[382] = 80'h8c1319;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[382] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[383] = 80'h725176;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[383] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[384] = 80'h56cec2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[384] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[385] = 80'h639a04;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[385] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[386] = 80'h5327e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[386] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[387] = 80'h1462c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[387] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[388] = 80'hd89f5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[388] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[389] = 80'h3902ae;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[389] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[390] = 80'ha2cbeb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[390] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[391] = 80'hf6681;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[391] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[392] = 80'h5dcafd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[392] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[393] = 80'h691152;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[393] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[394] = 80'h76bcf7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[394] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[395] = 80'h655333;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[395] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[396] = 80'h67c107;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[396] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[397] = 80'hbd651c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[397] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[398] = 80'hd88fbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[398] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[399] = 80'h3fa26a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[399] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[400] = 80'hbe3762;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[400] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[401] = 80'hee1fc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[401] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[402] = 80'hb30bdf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[402] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[403] = 80'h977fec;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[403] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[404] = 80'hf34eee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[404] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[405] = 80'h88c78e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[405] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[406] = 80'h50186a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[406] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[407] = 80'h22c496;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[407] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[408] = 80'h74ba14;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[408] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[409] = 80'h5fa922;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[409] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[410] = 80'h9f94e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[410] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[411] = 80'h66d9fb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[411] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[412] = 80'h10bb50;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[412] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[413] = 80'h139b8e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[413] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[414] = 80'h34094f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[414] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[415] = 80'hf852df;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[415] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[416] = 80'hb4b4a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[416] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[417] = 80'h7de478;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[417] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[418] = 80'h3db18f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[418] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[419] = 80'hd272a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[419] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[420] = 80'h8fb4b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[420] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[421] = 80'h39e1a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[421] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[422] = 80'hbcc07b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[422] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[423] = 80'hb2ab05;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[423] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[424] = 80'hf3b478;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[424] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[425] = 80'h9c9331;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[425] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[426] = 80'h570f8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[426] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[427] = 80'h92489c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[427] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[428] = 80'hd0fc4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[428] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[429] = 80'h2acd7b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[429] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[430] = 80'hab42dd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[430] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[431] = 80'he77e1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[431] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[432] = 80'h81a3c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[432] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[433] = 80'h6cf1fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[433] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[434] = 80'h34d05e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[434] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[435] = 80'h2b443d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[435] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[436] = 80'h97d73f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[436] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[437] = 80'h158478;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[437] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[438] = 80'he145aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[438] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[439] = 80'h1c385e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[439] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[440] = 80'hadbce3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[440] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[441] = 80'hd72c20;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[441] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[442] = 80'h5a3b1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[442] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[443] = 80'h5eaede;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[443] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[444] = 80'h651848;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[444] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[445] = 80'h977b39;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[445] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[446] = 80'h5cea8e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[446] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[447] = 80'h3b6c9a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[447] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[448] = 80'h492ee4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[448] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[449] = 80'h9a047c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[449] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[450] = 80'h608036;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[450] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[451] = 80'hcbe70e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[451] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[452] = 80'h1eb27a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[452] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[453] = 80'h751c3a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[453] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[454] = 80'h2b749f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[454] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[455] = 80'h7ab9cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[455] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[456] = 80'hdb74b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[456] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[457] = 80'h38ccf5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[457] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[458] = 80'hb81901;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[458] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[459] = 80'hdb6f8a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[459] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[460] = 80'hbdfaee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[460] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[461] = 80'hab9134;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[461] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[462] = 80'h6d74aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[462] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[463] = 80'hf71076;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[463] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[464] = 80'h579bdc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[464] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[465] = 80'hbbbd64;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[465] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[466] = 80'h83ae74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[466] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[467] = 80'hf8c1d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[467] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[468] = 80'hc8ed3e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[468] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[469] = 80'h2bf8dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[469] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[470] = 80'h16e5de;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[470] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[471] = 80'hb99492;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[471] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[472] = 80'h820b16;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[472] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[473] = 80'h8ae9cf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[473] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[474] = 80'hf6aad1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[474] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[475] = 80'hdef433;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[475] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[476] = 80'h60e02b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[476] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[477] = 80'hba10d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[477] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[478] = 80'h125ae0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[478] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[479] = 80'h75abca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[479] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[480] = 80'h7d0a37;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[480] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[481] = 80'h76c3eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[481] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[482] = 80'hee5867;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[482] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[483] = 80'ha63aa9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[483] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[484] = 80'h3bf1a7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[484] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[485] = 80'h41b00e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[485] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[486] = 80'h5dfcea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[486] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[487] = 80'h856939;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[487] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[488] = 80'h7fdd0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[488] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[489] = 80'hcac855;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[489] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[490] = 80'h82c86b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[490] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[491] = 80'h7d64e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[491] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[492] = 80'hc05790;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[492] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[493] = 80'h41b488;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[493] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[494] = 80'h19ef12;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[494] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[495] = 80'h89d14b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[495] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[496] = 80'hb42732;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[496] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[497] = 80'ha795fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[497] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[498] = 80'ha72e70;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[498] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[499] = 80'ha16e73;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[499] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[500] = 80'h80fe5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[500] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[501] = 80'hbdf1f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[501] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[502] = 80'h24e03d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[502] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[503] = 80'hcd8833;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[503] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[504] = 80'hd48427;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[504] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[505] = 80'h29413e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[505] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[506] = 80'h99f215;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[506] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[507] = 80'h43ea2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[507] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[508] = 80'hb05ed6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[508] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[509] = 80'h359c4e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[509] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[510] = 80'ha53a50;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[510] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[511] = 80'hba0217;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[511] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[512] = 80'ha7a8be;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[512] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[513] = 80'h117261;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[513] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[514] = 80'hba40b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[514] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[515] = 80'hd3778c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[515] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[516] = 80'h133300;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[516] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[517] = 80'h8026d0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[517] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[518] = 80'h3c2a96;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[518] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[519] = 80'haf2172;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[519] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[520] = 80'hf83e69;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[520] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[521] = 80'h2bae72;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[521] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[522] = 80'haaffe3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[522] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[523] = 80'he47a3a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[523] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[524] = 80'hecf185;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[524] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[525] = 80'h2ed0f5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[525] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[526] = 80'hd53425;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[526] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[527] = 80'hecfd2a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[527] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[528] = 80'hc133a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[528] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[529] = 80'hb51947;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[529] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[530] = 80'h1f5b10;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[530] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[531] = 80'h724175;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[531] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[532] = 80'h4a6946;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[532] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[533] = 80'hf4634a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[533] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[534] = 80'h74e5f6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[534] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[535] = 80'hb53980;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[535] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[536] = 80'hbbd32a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[536] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[537] = 80'h4beff2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[537] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[538] = 80'hc8358f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[538] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[539] = 80'hcb9cd4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[539] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[540] = 80'h5a3371;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[540] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[541] = 80'hb24300;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[541] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[542] = 80'h1fb996;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[542] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[543] = 80'hbd4f61;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[543] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[544] = 80'h8abbcd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[544] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[545] = 80'hb9b2c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[545] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[546] = 80'h638408;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[546] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[547] = 80'hd821e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[547] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[548] = 80'h694d89;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[548] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[549] = 80'hcc2430;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[549] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[550] = 80'hb3c95;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[550] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[551] = 80'h2c40c9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[551] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[552] = 80'hec7053;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[552] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[553] = 80'h8adfbd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[553] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[554] = 80'h15e421;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[554] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[555] = 80'hcd639d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[555] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[556] = 80'h6a5ec;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[556] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[557] = 80'h4837b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[557] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[558] = 80'h3c1296;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[558] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[559] = 80'h9854db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[559] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[560] = 80'he23953;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[560] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[561] = 80'h6e5f61;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[561] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[562] = 80'hb67704;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[562] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[563] = 80'hc188f5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[563] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[564] = 80'h9f0af0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[564] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[565] = 80'h13deba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[565] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[566] = 80'hd836a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[566] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[567] = 80'h378015;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[567] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[568] = 80'h6857c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[568] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[569] = 80'h920848;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[569] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[570] = 80'hdf91e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[570] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[571] = 80'h203539;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[571] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[572] = 80'he0e16e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[572] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[573] = 80'h518348;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[573] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[574] = 80'h29589f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[574] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[575] = 80'hd5eff5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[575] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[576] = 80'ha8909a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[576] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[577] = 80'hc6ccb7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[577] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[578] = 80'h8fd56d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[578] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[579] = 80'hbf7f6d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[579] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[580] = 80'h6a229b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[580] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[581] = 80'ha7dd84;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[581] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[582] = 80'h3d9854;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[582] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[583] = 80'h3c87c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[583] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[584] = 80'h588ad5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[584] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[585] = 80'heaaf14;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[585] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[586] = 80'h344bf2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[586] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[587] = 80'h3d9161;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[587] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[588] = 80'h415ce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[588] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[589] = 80'hb69cc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[589] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[590] = 80'hfe9312;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[590] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[591] = 80'h878cb6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[591] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[592] = 80'h38cf4e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[592] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[593] = 80'h76dcb4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[593] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[594] = 80'h702f85;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[594] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[595] = 80'hecdc20;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[595] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[596] = 80'h64eed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[596] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[597] = 80'h197ad7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[597] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[598] = 80'h860fe2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[598] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[599] = 80'haafcfa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[599] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[600] = 80'hb3fdf0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[600] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[601] = 80'h75513;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[601] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[602] = 80'h13141b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[602] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[603] = 80'hd07c80;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[603] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[604] = 80'h7023d5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[604] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[605] = 80'h88bbc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[605] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[606] = 80'h8bd1c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[606] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[607] = 80'hede0cc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[607] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[608] = 80'h11d1b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[608] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[609] = 80'hd0feb3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[609] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[610] = 80'hef7aab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[610] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[611] = 80'h929846;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[611] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[612] = 80'h87f8f5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[612] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[613] = 80'hf6d906;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[613] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[614] = 80'h301023;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[614] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[615] = 80'hc0367e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[615] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[616] = 80'hb5225;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[616] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[617] = 80'h1abda8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[617] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[618] = 80'hf76cf7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[618] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[619] = 80'h715672;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[619] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[620] = 80'h7a6132;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[620] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[621] = 80'h443d93;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[621] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[622] = 80'heb213b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[622] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[623] = 80'h4d47a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[623] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[624] = 80'ha05377;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[624] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[625] = 80'h6ac1b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[625] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[626] = 80'h7a773d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[626] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[627] = 80'he5e3a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[627] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[628] = 80'hc9746b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[628] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[629] = 80'h23a9d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[629] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[630] = 80'h4ec356;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[630] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[631] = 80'h75d68;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[631] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[632] = 80'h3f8eba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[632] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[633] = 80'h4d98e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[633] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[634] = 80'h98da92;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[634] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[635] = 80'hca02ef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[635] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[636] = 80'h924656;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[636] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[637] = 80'h4eb306;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[637] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[638] = 80'h33a608;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[638] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[639] = 80'h291e21;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[639] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[640] = 80'hc4dc56;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[640] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[641] = 80'h1b53a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[641] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[642] = 80'h9d22f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[642] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[643] = 80'h5a1b8f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[643] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[644] = 80'he01679;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[644] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[645] = 80'h44e0ed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[645] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[646] = 80'hc9bb74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[646] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[647] = 80'h5c1683;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[647] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[648] = 80'h5fbc9d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[648] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[649] = 80'hbc2b03;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[649] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[650] = 80'h44df86;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[650] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[651] = 80'hdadec5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[651] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[652] = 80'h2fa3c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[652] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[653] = 80'h795c0b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[653] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[654] = 80'hc6f84e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[654] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[655] = 80'hb16934;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[655] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[656] = 80'h9460ec;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[656] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[657] = 80'h961e88;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[657] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[658] = 80'hc93603;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[658] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[659] = 80'hf71bb0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[659] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[660] = 80'hb1611c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[660] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[661] = 80'hec7932;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[661] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[662] = 80'h43bb09;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[662] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[663] = 80'h40cb8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[663] = 80'h7ffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[664] = 80'h85d475;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[664] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[665] = 80'ha661a8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[665] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[666] = 80'hf38b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[666] = 80'hfffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[667] = 80'h986622;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[667] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[668] = 80'h72876e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[668] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[669] = 80'h26c981;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[669] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[670] = 80'hc3c23a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[670] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[671] = 80'h907259;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[671] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[672] = 80'h52165d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[672] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[673] = 80'h95fcd7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[673] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[674] = 80'h2dc5de;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[674] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[675] = 80'h3bd5a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[675] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[676] = 80'ha551ba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[676] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[677] = 80'h35e5cb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[677] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[678] = 80'hc960bd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[678] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[679] = 80'h23b8b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[679] = 80'h3fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[680] = 80'hd4d778;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[680] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[681] = 80'hea3ee3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[681] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[682] = 80'h1d84d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[682] = 80'h1fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[683] = 80'h77135c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[683] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[684] = 80'h61df00;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[684] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[685] = 80'ha9a5bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[685] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[686] = 80'hba4d19;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[686] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[687] = 80'hccf409;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[687] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[688] = 80'h85da8d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[688] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[689] = 80'h615d80;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[689] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[690] = 80'h726469;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[690] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[691] = 80'h69cc0a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[691] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[692] = 80'hb23db7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[692] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[693] = 80'h512c45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[693] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[694] = 80'hdcffc3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[694] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[695] = 80'hcc8fd4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[695] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[696] = 80'hac910e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[696] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[697] = 80'h66efed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[697] = 80'h7fffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[698] = 80'hd0094e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[698] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[699] = 80'hc23370;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[699] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem[700] = 80'hace597;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[5].u_tcam.mem_mask[700] = 80'hffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[1] = 80'hc76428a3ac18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[1] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[2] = 80'h6fa2b332a044;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[2] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[3] = 80'hdf160ea7e244;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[3] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[4] = 80'hbde8a5158a2b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[4] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[5] = 80'h1c7fcaa5772f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[5] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[6] = 80'h398bc2065413;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[6] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[7] = 80'hbf26a132d23e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[7] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[8] = 80'h2e5a52ddfb3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[8] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[9] = 80'hf9c4f448c4c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[9] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[10] = 80'h35e4dd182f90;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[10] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[11] = 80'h8513d0c50521;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[11] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[12] = 80'h35a66285b62e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[12] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[13] = 80'h4915d9de428f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[13] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[14] = 80'h3eff489073c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[14] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[15] = 80'hd00165db49c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[15] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[16] = 80'hc6e7d540048a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[16] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[17] = 80'hd2cf31221e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[17] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[18] = 80'h9cc2400c08bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[18] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[19] = 80'he84ab68b1a24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[19] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[20] = 80'hdc9c606e91ae;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[20] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[21] = 80'h4b8ee53f7660;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[21] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[22] = 80'ha6dc109cdbbd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[22] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[23] = 80'h2e5acd726cb2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[23] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[24] = 80'hbb30b2ecd487;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[24] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[25] = 80'h9aeec82f8fac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[25] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[26] = 80'hab83fe2b985c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[26] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[27] = 80'hca3daac02b2f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[27] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[28] = 80'h1a893b2ffa10;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[28] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[29] = 80'hcb1ab883d9ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[29] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[30] = 80'h6ddb0412e88d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[30] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[31] = 80'h25d034a677c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[31] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[32] = 80'h2ee63ce89af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[32] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[33] = 80'h1ab5a710d843;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[33] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[34] = 80'h97e8c062f084;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[34] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[35] = 80'h30a809743d4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[35] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[36] = 80'h22420da7f8f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[36] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[37] = 80'hafaf284ad3bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[37] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[38] = 80'h53bd4f0d7794;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[38] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[39] = 80'h5c0d39f2f061;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[39] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[40] = 80'h9419a7ce074a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[40] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[41] = 80'h52d45cc1e4a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[41] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[42] = 80'h9b30665b9971;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[42] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[43] = 80'h20d936f412c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[43] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[44] = 80'h8b889af41550;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[44] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[45] = 80'hf91ce85e797d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[45] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[46] = 80'h6e1dbd81191;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[46] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[47] = 80'h345e3c5f1365;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[47] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[48] = 80'h8dceefe91dc9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[48] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[49] = 80'hd47d2191ffed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[49] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[50] = 80'h7d341fbc821b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[50] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[51] = 80'h2e1c5d9ff7d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[51] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[52] = 80'hb7c667fd0324;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[52] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[53] = 80'h4933bf21a16c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[53] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[54] = 80'hf9724902347e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[54] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[55] = 80'haeb766b220db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[55] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[56] = 80'hdbbc2a3224ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[56] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[57] = 80'h365a679e8085;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[57] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[58] = 80'heeff7c2b7b33;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[58] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[59] = 80'h45bb6a31bb68;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[59] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[60] = 80'h1a81b1c43f91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[60] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[61] = 80'h1de0ad29184a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[61] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[62] = 80'h4eb9229cd415;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[62] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[63] = 80'h75c39cfd15db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[63] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[64] = 80'hbd7d9ddf726;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[64] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[65] = 80'h788ece7eed43;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[65] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[66] = 80'h689790000fff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[66] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[67] = 80'h30fca31cf96b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[67] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[68] = 80'h358975cc2823;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[68] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[69] = 80'h6b1cd921c79d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[69] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[70] = 80'h549a31ff63b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[70] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[71] = 80'h310dee607220;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[71] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[72] = 80'haf90fc2fb606;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[72] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[73] = 80'hdb655000d3a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[73] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[74] = 80'h8bf35344ab45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[74] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[75] = 80'h2d8a38190b20;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[75] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[76] = 80'h263f7f66582;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[76] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[77] = 80'h4dfc2ba4768d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[77] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[78] = 80'h849983bfbe7a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[78] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[79] = 80'h1efcb2f4dd4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[79] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[80] = 80'h61e5a9de4569;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[80] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[81] = 80'h770c1c4bd3a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[81] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[82] = 80'h500562660aff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[82] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[83] = 80'ha72a189143e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[83] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[84] = 80'h51a64abf0e09;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[84] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[85] = 80'h1f5700abe928;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[85] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[86] = 80'h512e72fad6a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[86] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[87] = 80'h5f3a530396cf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[87] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[88] = 80'h748487400445;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[88] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[89] = 80'h87719fb3f864;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[89] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[90] = 80'he88c8f60061d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[90] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[91] = 80'h9f6cc5f93019;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[91] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[92] = 80'hfa9df2c0fa11;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[92] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[93] = 80'h3e5de237f4f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[93] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[94] = 80'h1220e6f8b9fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[94] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[95] = 80'hceb0c2f94c3c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[95] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[96] = 80'h1845b8356ded;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[96] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[97] = 80'hcb7d6f052ed9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[97] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[98] = 80'ha1d827523dc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[98] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[99] = 80'hcaf8264a3ea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[99] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[100] = 80'h38ead3f12916;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[100] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[101] = 80'h13d2ee37c448;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[101] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[102] = 80'h3c2fe7d9f34c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[102] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[103] = 80'h3c1db8626079;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[103] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[104] = 80'h865b861ca607;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[104] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[105] = 80'h794600c6d0f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[105] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[106] = 80'he00c57f6e0b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[106] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[107] = 80'he29db65e8903;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[107] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[108] = 80'h8e261e6170f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[108] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[109] = 80'h66939b10ec73;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[109] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[110] = 80'h70c2e9c3c8eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[110] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[111] = 80'h45c66be84cf4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[111] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[112] = 80'h232cef211d0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[112] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[113] = 80'h80542dda5aa2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[113] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[114] = 80'h474effbc30dd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[114] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[115] = 80'he4cebd5c6fa4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[115] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[116] = 80'haf6a54830375;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[116] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[117] = 80'h8ef028be44c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[117] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[118] = 80'h5fdca8436bf4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[118] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[119] = 80'h6e7e1c15bd08;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[119] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[120] = 80'h134c1f65fd66;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[120] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[121] = 80'hcea87493679f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[121] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[122] = 80'hceb7bc309c1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[122] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[123] = 80'h61a6f8771878;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[123] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[124] = 80'hcedef6a567fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[124] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[125] = 80'h2e32a08622cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[125] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[126] = 80'h5356e16b8fd7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[126] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[127] = 80'hfd605bd942c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[127] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[128] = 80'hd5f103f449;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[128] = 80'hffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[129] = 80'h5f57f4362b22;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[129] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[130] = 80'h2e67f284f871;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[130] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[131] = 80'hecd79dcadc01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[131] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[132] = 80'he00525c7b0f8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[132] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[133] = 80'hb3cf483e6c80;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[133] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[134] = 80'h77eb26f31bbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[134] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[135] = 80'h8b676c49d915;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[135] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[136] = 80'ha2822acbd35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[136] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[137] = 80'h3a257929df1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[137] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[138] = 80'he9b0e1c40a18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[138] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[139] = 80'h3f10a0b32f42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[139] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[140] = 80'hf8a042a8b1d1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[140] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[141] = 80'hc010041f98fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[141] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[142] = 80'h6f5155d6bf2a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[142] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[143] = 80'h6174e0aee88e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[143] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[144] = 80'hd8f296505931;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[144] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[145] = 80'he512e3c64789;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[145] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[146] = 80'h373e0b9976b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[146] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[147] = 80'h3e7dacda18b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[147] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[148] = 80'h964ddbc00a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[148] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[149] = 80'h54781b947c65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[149] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[150] = 80'h4e476ae23070;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[150] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[151] = 80'h965a202c5dd1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[151] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[152] = 80'h6eeef25e5a0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[152] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[153] = 80'hbd9be825e53c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[153] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[154] = 80'h5a0d2b0e2652;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[154] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[155] = 80'hf02c2960a78f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[155] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[156] = 80'h43801573ed5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[156] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[157] = 80'h34d1a3628645;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[157] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[158] = 80'h476d2c7ebc16;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[158] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[159] = 80'ha17de6c9b9c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[159] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[160] = 80'h2e3b2da7cb0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[160] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[161] = 80'h618fe75b3a00;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[161] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[162] = 80'h7868e9b929a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[162] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[163] = 80'hcbe5e4137d1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[163] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[164] = 80'h6771e8c490b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[164] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[165] = 80'h7be9cc15dbad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[165] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[166] = 80'h8c89b097b14c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[166] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[167] = 80'hf2124342ae18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[167] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[168] = 80'h330261ba3670;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[168] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[169] = 80'h42c4edb6d896;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[169] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[170] = 80'h23a570bc32da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[170] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[171] = 80'hdb4f2973fc73;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[171] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[172] = 80'h4c40d88318b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[172] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[173] = 80'h1273739101e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[173] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[174] = 80'h9c2ebac8770d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[174] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[175] = 80'haaeaffde1744;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[175] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[176] = 80'h67b1d0406ac4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[176] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[177] = 80'h602be7c25423;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[177] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[178] = 80'h7bd2374d89da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[178] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[179] = 80'h484efbf68ee5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[179] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[180] = 80'h8c2970d5df55;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[180] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[181] = 80'haec65cebfe7b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[181] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[182] = 80'h94dfc4cad63a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[182] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[183] = 80'h16398c9c5329;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[183] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[184] = 80'hc1d9c5b84501;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[184] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[185] = 80'hd1ad3332662b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[185] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[186] = 80'hb91d094ca5fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[186] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[187] = 80'h66807169ce5b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[187] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[188] = 80'h6ef096e4f564;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[188] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[189] = 80'h328864e675f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[189] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[190] = 80'h7dae2b0e1b45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[190] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[191] = 80'hbcb94b47b6e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[191] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[192] = 80'h969630df4be5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[192] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[193] = 80'h8fa1021a531a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[193] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[194] = 80'h872d61d5debf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[194] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[195] = 80'h991610788933;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[195] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[196] = 80'habf899e0a35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[196] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[197] = 80'h9a50b37b4c4e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[197] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[198] = 80'ha57859f9c477;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[198] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[199] = 80'h79cd60c49c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[199] = 80'h7fffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[200] = 80'h116a5a1abd7d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[200] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[201] = 80'hc21fd0b46818;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[201] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[202] = 80'hcb7c1d8cfffa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[202] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[203] = 80'h5da2668e789f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[203] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[204] = 80'ha975554d1660;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[204] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[205] = 80'hf527f8412a24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[205] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[206] = 80'h6e7cabe12a47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[206] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[207] = 80'hecce1c4cd86e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[207] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[208] = 80'h72d3d3fcd72b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[208] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[209] = 80'h839e1fb55d44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[209] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[210] = 80'h478398e0b9ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[210] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[211] = 80'h8530d50e759f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[211] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[212] = 80'h11f968361ebd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[212] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[213] = 80'h8ce994cc083f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[213] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[214] = 80'h2c23f84988ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[214] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[215] = 80'h9760938f25c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[215] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[216] = 80'h274efbfa8211;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[216] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[217] = 80'h694132b93ba3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[217] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[218] = 80'h682f3056401;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[218] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[219] = 80'hd1c36a785d4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[219] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[220] = 80'h4ae9b6d2ef4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[220] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[221] = 80'hc9c32ab41eeb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[221] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[222] = 80'hcbc076ebe28e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[222] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[223] = 80'hfbda31fd76c0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[223] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[224] = 80'h9a099a151b35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[224] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[225] = 80'h54a1681b3ffb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[225] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[226] = 80'hf0cf8f9ee272;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[226] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[227] = 80'h3f535b44d28a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[227] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[228] = 80'h7ae44fa333c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[228] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[229] = 80'hb665ce7f735a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[229] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[230] = 80'h626c7ae8774d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[230] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[231] = 80'hf3cddb51d392;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[231] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[232] = 80'h944a75a8319c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[232] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[233] = 80'heaacb9890fae;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[233] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[234] = 80'h46f6540ec7f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[234] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[235] = 80'hc6088fc1bd3d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[235] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[236] = 80'h5e0b61c56031;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[236] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[237] = 80'h27b4c51c3bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[237] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[238] = 80'hbe4d82d7e60e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[238] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[239] = 80'h7eef6a0932c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[239] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[240] = 80'h564f40cb3bc6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[240] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[241] = 80'h49ba0e14ede1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[241] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[242] = 80'hffa1385e8e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[242] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[243] = 80'hc2a6a6c5875c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[243] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[244] = 80'h46ed88992ff9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[244] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[245] = 80'h7bd52c488741;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[245] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[246] = 80'hdd037b320186;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[246] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[247] = 80'hbc45bae8ac0a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[247] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[248] = 80'h5b06c7e96f30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[248] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[249] = 80'hd4ddc557a673;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[249] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[250] = 80'h53ec21af6aa7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[250] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[251] = 80'h17ac57f88e87;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[251] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[252] = 80'ha4100e4032cc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[252] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[253] = 80'h140fa51dda60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[253] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[254] = 80'hba76b63b04af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[254] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[255] = 80'h7bf30212d42d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[255] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[256] = 80'h389a856d0929;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[256] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[257] = 80'h971def77bfa0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[257] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[258] = 80'h7fea6ca2dda9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[258] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[259] = 80'h6cc87b7163e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[259] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[260] = 80'h652f37432033;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[260] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[261] = 80'h94ca0afeaf40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[261] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[262] = 80'haa6075a82cfd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[262] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[263] = 80'he393132fbd4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[263] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[264] = 80'h8617fb8769a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[264] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[265] = 80'hd45704f554fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[265] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[266] = 80'h83aeac67707;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[266] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[267] = 80'had11dd592c9a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[267] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[268] = 80'h199fcd09ed28;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[268] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[269] = 80'h306fc67d4fd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[269] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[270] = 80'hded308236673;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[270] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[271] = 80'h6bb4f3981543;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[271] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[272] = 80'h28d774fa8bab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[272] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[273] = 80'h5f39e126fa40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[273] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[274] = 80'h4ec1930dd830;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[274] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[275] = 80'h2eabafa47444;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[275] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[276] = 80'hf2c4354979b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[276] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[277] = 80'h4375ff2839ff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[277] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[278] = 80'h831847d750e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[278] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[279] = 80'h6d4ff70a7fc3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[279] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[280] = 80'h67633ad96690;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[280] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[281] = 80'h58b1bb7ab35b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[281] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[282] = 80'h378d65b1297a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[282] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[283] = 80'h8ab24a720a34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[283] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[284] = 80'h9b617faf808a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[284] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[285] = 80'h2b5be33345f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[285] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[286] = 80'h80b069925240;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[286] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[287] = 80'h64819ae5ce38;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[287] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[288] = 80'hc8a2886319ad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[288] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[289] = 80'hbba80680cd74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[289] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[290] = 80'hc624c1780420;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[290] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[291] = 80'hdf4dc19f8a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[291] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[292] = 80'hbf4fc4c5109d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[292] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[293] = 80'h230e53a6e40d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[293] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[294] = 80'h6a8845704812;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[294] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[295] = 80'hd02d7e61c3ff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[295] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[296] = 80'h42d9ad4b7cb5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[296] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[297] = 80'h6620c43e40cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[297] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[298] = 80'h572b2a5075a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[298] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[299] = 80'hbc0a3cd8632;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[299] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[300] = 80'h318840f45c23;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[300] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[301] = 80'h7ec0b9f2df84;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[301] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[302] = 80'h708eaeea371;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[302] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[303] = 80'h29e3e9901c1f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[303] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[304] = 80'hf4f0fb40376f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[304] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[305] = 80'h7de8c27c7bf8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[305] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[306] = 80'h722214538bb3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[306] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[307] = 80'hb35284a2e8f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[307] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[308] = 80'hc1e963dc4088;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[308] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[309] = 80'h50d5503770e6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[309] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[310] = 80'hb63951662a30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[310] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[311] = 80'h7eddea567619;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[311] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[312] = 80'h4eab0a109e8f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[312] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[313] = 80'he549f26a551a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[313] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[314] = 80'h161e12d7d5f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[314] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[315] = 80'h2fb8691cf03d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[315] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[316] = 80'h6d0dd414bd88;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[316] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[317] = 80'hd47f0cfd8269;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[317] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[318] = 80'he7fe58f76aac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[318] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[319] = 80'hcddb5437e4b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[319] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[320] = 80'h58ac2d7d65c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[320] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[321] = 80'he81d8eb85034;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[321] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[322] = 80'ha6fb99d69d1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[322] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[323] = 80'h85db0f2ad52e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[323] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[324] = 80'hba447f49c0b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[324] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[325] = 80'h99d3496acd35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[325] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[326] = 80'h40e7e1b07303;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[326] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[327] = 80'h55f948ebe91d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[327] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[328] = 80'h392c0459ce02;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[328] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[329] = 80'h7e3d419f5d34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[329] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[330] = 80'he74efb58eaa7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[330] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[331] = 80'hf83f581e4482;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[331] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[332] = 80'h9cce1dfeef14;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[332] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[333] = 80'h4b70936e9f64;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[333] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[334] = 80'h8f60bf446783;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[334] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[335] = 80'h93a9046448e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[335] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[336] = 80'h6e3ce4ac6730;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[336] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[337] = 80'h84de22fbc40a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[337] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[338] = 80'h2d98732c0914;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[338] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[339] = 80'h588e0584287c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[339] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[340] = 80'h8f50e0497e89;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[340] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[341] = 80'hb0e119fb2555;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[341] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[342] = 80'h4cd3c2cde21a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[342] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[343] = 80'hda342cb3beee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[343] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[344] = 80'h9f7fc5e6a042;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[344] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[345] = 80'hcc5300c82669;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[345] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[346] = 80'h6a1ec386bf00;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[346] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[347] = 80'h2317e8d90545;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[347] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[348] = 80'h8d4fe98625cf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[348] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[349] = 80'h60665e2c19e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[349] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[350] = 80'h596674fbbfb1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[350] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[351] = 80'h5c7688d8aad5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[351] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[352] = 80'h99c3cb202d30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[352] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[353] = 80'ha86ac83a7681;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[353] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[354] = 80'hf9f330aaf7e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[354] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[355] = 80'h3c3dcdb988e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[355] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[356] = 80'h82440e73e0a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[356] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[357] = 80'hdeb63d376bdd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[357] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[358] = 80'h3f13c6d986da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[358] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[359] = 80'h959a11161a8a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[359] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[360] = 80'h4fc4b9709a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[360] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[361] = 80'h603260a4fa8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[361] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[362] = 80'h317642426d30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[362] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[363] = 80'h93eea5159da0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[363] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[364] = 80'ha6a6c5effbb8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[364] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[365] = 80'h9a556fc0f1e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[365] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[366] = 80'hca8bfde422b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[366] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[367] = 80'h6b3d4da4a0e4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[367] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[368] = 80'hb8725432eee0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[368] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[369] = 80'h2a5f4d97572c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[369] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[370] = 80'h3f4b2f37c91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[370] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[371] = 80'h6d012a56f306;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[371] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[372] = 80'hf39c18ff7423;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[372] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[373] = 80'h64fe54c3d020;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[373] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[374] = 80'h5941386df853;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[374] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[375] = 80'hfd5081a7023d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[375] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[376] = 80'h59d252677e44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[376] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[377] = 80'hb1ef710456c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[377] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[378] = 80'h8a3b29afa55f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[378] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[379] = 80'ha8f4af7c920a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[379] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[380] = 80'h9b5b556528f0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[380] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[381] = 80'h8d75c4ce6384;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[381] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[382] = 80'h644e172a4d39;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[382] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[383] = 80'h4e2c31c4e9bf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[383] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[384] = 80'hfb16e104670e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[384] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[385] = 80'hedda66338267;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[385] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[386] = 80'h28c12a16f1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[386] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[387] = 80'hff84824ad314;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[387] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[388] = 80'hbe7756aeeab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[388] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[389] = 80'h7e61e055303f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[389] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[390] = 80'haac7193a22af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[390] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[391] = 80'h565f0106873e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[391] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[392] = 80'h75032e61802d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[392] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[393] = 80'hf2f7c9dbbf6e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[393] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[394] = 80'hc616b82074dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[394] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[395] = 80'h9b90c73a26b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[395] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[396] = 80'hf1aad48501e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[396] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[397] = 80'hb50e5a5b2331;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[397] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[398] = 80'h536e70ff511;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[398] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[399] = 80'h500f137223d6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[399] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[400] = 80'h2791051b62a6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[400] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[401] = 80'hc4eb2c045df0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[401] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[402] = 80'ha4ad1b4e4c65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[402] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[403] = 80'h5dcd203c62ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[403] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[404] = 80'hbd2053fe1aa1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[404] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[405] = 80'hdd873733eebd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[405] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[406] = 80'hd5cc8944cc44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[406] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[407] = 80'hdf75e34c1d60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[407] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[408] = 80'h69516c90e02b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[408] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[409] = 80'hba7434218648;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[409] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[410] = 80'h75995e082cc9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[410] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[411] = 80'h8f8a0618c492;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[411] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[412] = 80'h85652adefb50;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[412] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[413] = 80'h84e3bbb346a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[413] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[414] = 80'hce288545ff5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[414] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[415] = 80'hf34840529bc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[415] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[416] = 80'h93b680734ca8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[416] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[417] = 80'h6d3e5930bf31;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[417] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[418] = 80'h4c6bb4e13dd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[418] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[419] = 80'hc17e7cae146d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[419] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[420] = 80'h3a01e234f448;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[420] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[421] = 80'h1f6089a70d31;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[421] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[422] = 80'he9910acedf01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[422] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[423] = 80'h92c1be63a45c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[423] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[424] = 80'h77250b5545e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[424] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[425] = 80'h41875a4af1b4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[425] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[426] = 80'h1f7188b8f195;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[426] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[427] = 80'he7043697f5e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[427] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[428] = 80'hccb0a5325cbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[428] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[429] = 80'hf77c99d0ae10;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[429] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[430] = 80'h51c66267cec7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[430] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[431] = 80'ha3eb7b517f7d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[431] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[432] = 80'h5e4b84a9a324;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[432] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[433] = 80'h263366d9a934;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[433] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[434] = 80'h35cd167e2bad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[434] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[435] = 80'hb2c3bbf8fba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[435] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[436] = 80'h8f19a66976c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[436] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[437] = 80'he0b42c35622b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[437] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[438] = 80'hdca9a6f1782c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[438] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[439] = 80'h9a1541c274a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[439] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[440] = 80'h44768a38b95d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[440] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[441] = 80'h38f48a68b142;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[441] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[442] = 80'h9759c188b4fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[442] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[443] = 80'ha08c0f3399b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[443] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[444] = 80'h820dea118ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[444] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[445] = 80'h786f4fec3569;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[445] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[446] = 80'h35502a9bf339;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[446] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[447] = 80'hede032f81911;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[447] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[448] = 80'h5d2da41d57;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[448] = 80'h7fffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[449] = 80'h1d551e45233a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[449] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[450] = 80'h1232e7e21619;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[450] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[451] = 80'h9656bf8e0b9d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[451] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[452] = 80'h282df63c9a42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[452] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[453] = 80'hfb8cfa3efc1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[453] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[454] = 80'he202a5e04142;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[454] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[455] = 80'hce14bd93ed55;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[455] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[456] = 80'hb29b6b75332;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[456] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[457] = 80'ha560cfe7acfc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[457] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[458] = 80'h99c7f0448e01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[458] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[459] = 80'h1dc007e9c85a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[459] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[460] = 80'hd5bbfcebded1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[460] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[461] = 80'h7a59ce859cc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[461] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[462] = 80'h4ea8c5b70bda;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[462] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[463] = 80'h52f1807fc08a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[463] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[464] = 80'h206171d9529a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[464] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[465] = 80'h498a7ea9d6a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[465] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[466] = 80'h68b1d8990008;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[466] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[467] = 80'hdfdd7f5c6649;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[467] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[468] = 80'h423c83f43d47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[468] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[469] = 80'h71daa74440c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[469] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[470] = 80'h6b7caeb2cb69;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[470] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[471] = 80'h9301716b199f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[471] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[472] = 80'hf30c2c261355;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[472] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[473] = 80'he1037b5789b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[473] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[474] = 80'h4ac85c163c30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[474] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[475] = 80'hbd2e17a3bd71;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[475] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[476] = 80'h8cfbaac12a25;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[476] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[477] = 80'he07f86b355a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[477] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[478] = 80'he24b3b5f435d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[478] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[479] = 80'hc6100a3221e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[479] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[480] = 80'hd601e9e5d6ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[480] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[481] = 80'ha2ee82f9007b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[481] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[482] = 80'hb4baf8944204;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[482] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[483] = 80'h78c5ee1f506d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[483] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[484] = 80'h94176a64d950;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[484] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[485] = 80'hbdc7edf2bed3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[485] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[486] = 80'hf6141087125a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[486] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[487] = 80'h4d8a6c4bb175;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[487] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[488] = 80'hd702b7ff755e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[488] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[489] = 80'h17ad459c4491;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[489] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[490] = 80'hbecd69de0af5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[490] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[491] = 80'h6db83a09cb40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[491] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[492] = 80'hc15a3192c54e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[492] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[493] = 80'h372729de79a7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[493] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[494] = 80'hb7d5a573112e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[494] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[495] = 80'he7598a8d64ef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[495] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[496] = 80'h4d77a8f186e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[496] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[497] = 80'hb3a7e8c62438;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[497] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[498] = 80'h5e628e40bad8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[498] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[499] = 80'h2c6ae9566a81;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[499] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[500] = 80'h7c8088a4d780;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[500] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[501] = 80'h449da718991b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[501] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[502] = 80'heb14915c851e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[502] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[503] = 80'h3527b3d245b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[503] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[504] = 80'h85d7cc131a8a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[504] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[505] = 80'hb448dcc734b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[505] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[506] = 80'h463282aaf56;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[506] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[507] = 80'he6f6fe35b667;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[507] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[508] = 80'h80c258b15826;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[508] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[509] = 80'hfaac4f7283f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[509] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[510] = 80'ha03cce697a88;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[510] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[511] = 80'hdf03c7e186d0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[511] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[512] = 80'hc301b2ddb491;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[512] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[513] = 80'h5a553a6d946;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[513] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[514] = 80'hec81a0ecf565;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[514] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[515] = 80'h25b7ba6c7a22;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[515] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[516] = 80'hff62f77af68e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[516] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[517] = 80'h90696c0e7c49;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[517] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[518] = 80'hdb542752b51b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[518] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[519] = 80'h5c669d7e5719;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[519] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[520] = 80'h7869b90d6d6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[520] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[521] = 80'h6ab3f4028bc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[521] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[522] = 80'hfaf254c81784;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[522] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[523] = 80'he91e80ddf2b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[523] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[524] = 80'h12ec8002dccf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[524] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[525] = 80'h1fb66119b301;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[525] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[526] = 80'h35cfa56dca6a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[526] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[527] = 80'h257f17287640;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[527] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[528] = 80'he24b719e5fd5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[528] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[529] = 80'h1b6de98d63bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[529] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[530] = 80'hc7396a1e1d0b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[530] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[531] = 80'h7fb43ae9cd4b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[531] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[532] = 80'ha389a8825008;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[532] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[533] = 80'h62002cc089d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[533] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[534] = 80'ha2fc3e097fd8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[534] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[535] = 80'h93938f2e7bb6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[535] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[536] = 80'h4c0878c8f3c9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[536] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[537] = 80'h6dad4681d74b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[537] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[538] = 80'h90d849afd440;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[538] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[539] = 80'h99cea5c192b2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[539] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[540] = 80'h439a63924ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[540] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[541] = 80'h22efe4c3db4e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[541] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[542] = 80'h935f8ae1eaca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[542] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[543] = 80'h980ce89cb3ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[543] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[544] = 80'hb2b1d54e6143;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[544] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[545] = 80'h985262ca09c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[545] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[546] = 80'h1b5370c23148;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[546] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[547] = 80'hfa6e44897737;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[547] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[548] = 80'hedc347b5f551;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[548] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[549] = 80'hbbafbcb86844;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[549] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[550] = 80'h7fb9ba95cb59;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[550] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[551] = 80'hbe931b35ee21;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[551] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[552] = 80'h39f56d709e34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[552] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[553] = 80'h4e9dfa08200a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[553] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[554] = 80'h820c31b21a45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[554] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[555] = 80'h5c7809f7005;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[555] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[556] = 80'h3aca0c094cca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[556] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[557] = 80'h745ae42f60b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[557] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[558] = 80'h9ab1034e7c6e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[558] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[559] = 80'h8b03e00b02c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[559] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[560] = 80'h291393c268aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[560] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[561] = 80'h4f5dda910b46;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[561] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[562] = 80'hd702572b740;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[562] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[563] = 80'h82eb751a50eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[563] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[564] = 80'h69f1bf212be5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[564] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[565] = 80'h692f8eeae2e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[565] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[566] = 80'h19a683169415;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[566] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[567] = 80'h93bac3e6e685;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[567] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[568] = 80'h4993bee769ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[568] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[569] = 80'hcd7fb4cb6753;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[569] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[570] = 80'h240e7a3c36d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[570] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[571] = 80'hdee7cb29be85;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[571] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[572] = 80'h992597565e42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[572] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[573] = 80'h5cf48819c736;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[573] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[574] = 80'h47abe210da7f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[574] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[575] = 80'hf93a1757baa0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[575] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[576] = 80'h7c1ceb4afc56;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[576] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[577] = 80'haf7d256d7cc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[577] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[578] = 80'h56f4eacb32c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[578] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[579] = 80'hb0d1add53e47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[579] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[580] = 80'hd2755cc4bd17;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[580] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[581] = 80'ha6985589f9f2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[581] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[582] = 80'hc617a79d7ece;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[582] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[583] = 80'hce74602fffba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[583] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[584] = 80'hf924b4b96d61;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[584] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[585] = 80'h8c0b6b9901dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[585] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[586] = 80'hf68af87708bf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[586] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[587] = 80'h74fa5f30fe3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[587] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[588] = 80'h4db8a921b1d2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[588] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[589] = 80'h18a72f979e24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[589] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[590] = 80'h595e18260e26;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[590] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[591] = 80'haad2d483e822;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[591] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[592] = 80'h343913fad305;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[592] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[593] = 80'hb3d2b6c10e97;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[593] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[594] = 80'h5b359f4f70b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[594] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[595] = 80'h910fdf65238e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[595] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[596] = 80'h858d2a03d342;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[596] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[597] = 80'h60c0b6079327;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[597] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[598] = 80'hac7bf03559d7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[598] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[599] = 80'h9ad2390bbe32;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[599] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[600] = 80'hfa4f7ce06718;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[600] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[601] = 80'hd16fe65ec39f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[601] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[602] = 80'h2d99e55053a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[602] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[603] = 80'h5159029f3697;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[603] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[604] = 80'hb4b0447b5549;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[604] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[605] = 80'h377b752a37b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[605] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[606] = 80'h220bb11437f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[606] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[607] = 80'habd69fb1204e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[607] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[608] = 80'heb47988d0d8b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[608] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[609] = 80'hca9cc767edce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[609] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[610] = 80'h3b6f42cbe0a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[610] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[611] = 80'h1dd3fa287076;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[611] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[612] = 80'h9628912dbff2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[612] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[613] = 80'h89a7951bea35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[613] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[614] = 80'hc7b2ff90ab75;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[614] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[615] = 80'h7ec37d3f35d1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[615] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[616] = 80'h486d45350ba4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[616] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[617] = 80'hf7c78a4aeffd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[617] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[618] = 80'hea7f3c4470a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[618] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[619] = 80'h95398bca46db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[619] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[620] = 80'h2a21d269ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[620] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[621] = 80'h5ff142432afa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[621] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[622] = 80'h8d346fc65e2b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[622] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[623] = 80'h1a6584f50556;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[623] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[624] = 80'h8386da1029f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[624] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[625] = 80'hdb56c981ece6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[625] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[626] = 80'hcfe8af38f522;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[626] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[627] = 80'h8e919d8a745b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[627] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[628] = 80'h543818958c78;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[628] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[629] = 80'ha8b931f97188;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[629] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[630] = 80'h7dee0d849922;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[630] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[631] = 80'h1017ca8a2953;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[631] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[632] = 80'h7ed9cae24403;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[632] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[633] = 80'hea187ed4d55a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[633] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[634] = 80'h2e76e28270f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[634] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[635] = 80'hf1980343333f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[635] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[636] = 80'h8de1c963c062;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[636] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[637] = 80'h3fd86ea44501;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[637] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[638] = 80'hdc791a00bf2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[638] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[639] = 80'h76fd772b3105;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[639] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[640] = 80'h9137a6d429b2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[640] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[641] = 80'h49d4cbef7ccc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[641] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[642] = 80'h8051f12b529f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[642] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[643] = 80'h8d6aa657a5e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[643] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[644] = 80'h44bafb829ee6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[644] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[645] = 80'he55061ccc7b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[645] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[646] = 80'hd75970bd3bb0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[646] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[647] = 80'h4811729ba385;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[647] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[648] = 80'hc0501fd955df;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[648] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[649] = 80'h659c29b06d69;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[649] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[650] = 80'h6aec373261a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[650] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[651] = 80'hc25cd90f5dab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[651] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[652] = 80'hcee3230bfef6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[652] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[653] = 80'h7bde198a992f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[653] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[654] = 80'h7cd4d9587ccb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[654] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[655] = 80'h5cee7e94dd42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[655] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[656] = 80'hc7f2c96b613;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[656] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[657] = 80'hf2de9d0bdde4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[657] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[658] = 80'hb80342294761;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[658] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[659] = 80'hef05f9051dde;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[659] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[660] = 80'h89d9864b0f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[660] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[661] = 80'hf84ebc6b5933;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[661] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[662] = 80'h99c7ebd6ef11;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[662] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[663] = 80'ha5cfc726453c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[663] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[664] = 80'h8e33ccc43905;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[664] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[665] = 80'h61dbc393f8b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[665] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[666] = 80'hb5776eb8e40c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[666] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[667] = 80'hc56f02fbb8af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[667] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[668] = 80'hf06ac89a6e2e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[668] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[669] = 80'h4d46ea5704c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[669] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[670] = 80'h18a0d2ab536;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[670] = 80'h1ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[671] = 80'hde24ea9c8559;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[671] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[672] = 80'h117c2dcb8a3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[672] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[673] = 80'h42c5800a198;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[673] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[674] = 80'hc866641162c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[674] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[675] = 80'hc59ce2a178ef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[675] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[676] = 80'h91b9a88b2186;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[676] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[677] = 80'hbaaaa92f9330;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[677] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[678] = 80'h899bc4d45fed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[678] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[679] = 80'h31aba86c07cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[679] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[680] = 80'hc4984e56b9a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[680] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[681] = 80'h1b2cb5378bd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[681] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[682] = 80'hff120ca68f9a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[682] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[683] = 80'ha835dfd4a64e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[683] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[684] = 80'hcc35683c57dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[684] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[685] = 80'ha5c1099a0ccc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[685] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[686] = 80'hefd95c4e5fe9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[686] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[687] = 80'h7c76d25796aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[687] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[688] = 80'h7b60730923d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[688] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[689] = 80'h7373b8b8f3c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[689] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[690] = 80'h37e56c799b77;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[690] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[691] = 80'h64aeec7ab84c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[691] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[692] = 80'hdc1814387312;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[692] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[693] = 80'hdd2835b8c4f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[693] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[694] = 80'h5af2eb552cca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[694] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[695] = 80'h446b9299fa74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[695] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[696] = 80'h86928cf64fc6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[696] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[697] = 80'hc4fdc019c61f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[697] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[698] = 80'h882f97bb161f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[698] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[699] = 80'h4ed606f4518d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[699] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem[700] = 80'hbd46a3aa3c15;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[6].u_tcam.mem_mask[700] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[1] = 80'hc76428a3ac18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[1] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[2] = 80'h6fa2b332a044;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[2] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[3] = 80'hdf160ea7e244;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[3] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[4] = 80'hbde8a5158a2b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[4] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[5] = 80'h1c7fcaa5772f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[5] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[6] = 80'h398bc2065413;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[6] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[7] = 80'hbf26a132d23e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[7] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[8] = 80'h2e5a52ddfb3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[8] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[9] = 80'hf9c4f448c4c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[9] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[10] = 80'h35e4dd182f90;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[10] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[11] = 80'h8513d0c50521;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[11] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[12] = 80'h35a66285b62e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[12] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[13] = 80'h4915d9de428f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[13] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[14] = 80'h3eff489073c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[14] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[15] = 80'hd00165db49c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[15] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[16] = 80'hc6e7d540048a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[16] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[17] = 80'hd2cf31221e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[17] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[18] = 80'h9cc2400c08bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[18] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[19] = 80'he84ab68b1a24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[19] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[20] = 80'hdc9c606e91ae;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[20] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[21] = 80'h4b8ee53f7660;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[21] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[22] = 80'ha6dc109cdbbd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[22] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[23] = 80'h2e5acd726cb2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[23] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[24] = 80'hbb30b2ecd487;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[24] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[25] = 80'h9aeec82f8fac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[25] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[26] = 80'hab83fe2b985c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[26] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[27] = 80'hca3daac02b2f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[27] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[28] = 80'h1a893b2ffa10;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[28] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[29] = 80'hcb1ab883d9ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[29] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[30] = 80'h6ddb0412e88d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[30] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[31] = 80'h25d034a677c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[31] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[32] = 80'h2ee63ce89af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[32] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[33] = 80'h1ab5a710d843;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[33] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[34] = 80'h97e8c062f084;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[34] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[35] = 80'h30a809743d4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[35] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[36] = 80'h22420da7f8f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[36] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[37] = 80'hafaf284ad3bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[37] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[38] = 80'h53bd4f0d7794;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[38] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[39] = 80'h5c0d39f2f061;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[39] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[40] = 80'h9419a7ce074a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[40] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[41] = 80'h52d45cc1e4a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[41] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[42] = 80'h9b30665b9971;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[42] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[43] = 80'h20d936f412c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[43] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[44] = 80'h8b889af41550;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[44] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[45] = 80'hf91ce85e797d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[45] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[46] = 80'h6e1dbd81191;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[46] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[47] = 80'h345e3c5f1365;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[47] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[48] = 80'h8dceefe91dc9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[48] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[49] = 80'hd47d2191ffed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[49] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[50] = 80'h7d341fbc821b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[50] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[51] = 80'h2e1c5d9ff7d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[51] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[52] = 80'hb7c667fd0324;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[52] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[53] = 80'h4933bf21a16c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[53] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[54] = 80'hf9724902347e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[54] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[55] = 80'haeb766b220db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[55] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[56] = 80'hdbbc2a3224ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[56] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[57] = 80'h365a679e8085;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[57] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[58] = 80'heeff7c2b7b33;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[58] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[59] = 80'h45bb6a31bb68;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[59] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[60] = 80'h1a81b1c43f91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[60] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[61] = 80'h1de0ad29184a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[61] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[62] = 80'h4eb9229cd415;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[62] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[63] = 80'h75c39cfd15db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[63] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[64] = 80'hbd7d9ddf726;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[64] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[65] = 80'h788ece7eed43;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[65] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[66] = 80'h689790000fff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[66] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[67] = 80'h30fca31cf96b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[67] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[68] = 80'h358975cc2823;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[68] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[69] = 80'h6b1cd921c79d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[69] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[70] = 80'h549a31ff63b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[70] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[71] = 80'h310dee607220;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[71] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[72] = 80'haf90fc2fb606;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[72] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[73] = 80'hdb655000d3a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[73] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[74] = 80'h8bf35344ab45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[74] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[75] = 80'h2d8a38190b20;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[75] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[76] = 80'h263f7f66582;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[76] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[77] = 80'h4dfc2ba4768d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[77] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[78] = 80'h849983bfbe7a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[78] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[79] = 80'h1efcb2f4dd4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[79] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[80] = 80'h61e5a9de4569;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[80] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[81] = 80'h770c1c4bd3a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[81] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[82] = 80'h500562660aff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[82] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[83] = 80'ha72a189143e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[83] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[84] = 80'h51a64abf0e09;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[84] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[85] = 80'h1f5700abe928;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[85] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[86] = 80'h512e72fad6a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[86] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[87] = 80'h5f3a530396cf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[87] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[88] = 80'h748487400445;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[88] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[89] = 80'h87719fb3f864;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[89] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[90] = 80'he88c8f60061d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[90] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[91] = 80'h9f6cc5f93019;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[91] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[92] = 80'hfa9df2c0fa11;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[92] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[93] = 80'h3e5de237f4f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[93] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[94] = 80'h1220e6f8b9fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[94] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[95] = 80'hceb0c2f94c3c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[95] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[96] = 80'h1845b8356ded;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[96] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[97] = 80'hcb7d6f052ed9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[97] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[98] = 80'ha1d827523dc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[98] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[99] = 80'hcaf8264a3ea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[99] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[100] = 80'h38ead3f12916;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[100] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[101] = 80'h13d2ee37c448;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[101] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[102] = 80'h3c2fe7d9f34c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[102] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[103] = 80'h3c1db8626079;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[103] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[104] = 80'h865b861ca607;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[104] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[105] = 80'h794600c6d0f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[105] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[106] = 80'he00c57f6e0b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[106] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[107] = 80'he29db65e8903;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[107] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[108] = 80'h8e261e6170f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[108] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[109] = 80'h66939b10ec73;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[109] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[110] = 80'h70c2e9c3c8eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[110] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[111] = 80'h45c66be84cf4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[111] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[112] = 80'h232cef211d0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[112] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[113] = 80'h80542dda5aa2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[113] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[114] = 80'h474effbc30dd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[114] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[115] = 80'he4cebd5c6fa4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[115] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[116] = 80'haf6a54830375;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[116] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[117] = 80'h8ef028be44c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[117] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[118] = 80'h5fdca8436bf4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[118] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[119] = 80'h6e7e1c15bd08;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[119] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[120] = 80'h134c1f65fd66;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[120] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[121] = 80'hcea87493679f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[121] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[122] = 80'hceb7bc309c1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[122] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[123] = 80'h61a6f8771878;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[123] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[124] = 80'hcedef6a567fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[124] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[125] = 80'h2e32a08622cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[125] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[126] = 80'h5356e16b8fd7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[126] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[127] = 80'hfd605bd942c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[127] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[128] = 80'hd5f103f449;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[128] = 80'hffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[129] = 80'h5f57f4362b22;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[129] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[130] = 80'h2e67f284f871;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[130] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[131] = 80'hecd79dcadc01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[131] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[132] = 80'he00525c7b0f8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[132] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[133] = 80'hb3cf483e6c80;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[133] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[134] = 80'h77eb26f31bbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[134] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[135] = 80'h8b676c49d915;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[135] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[136] = 80'ha2822acbd35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[136] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[137] = 80'h3a257929df1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[137] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[138] = 80'he9b0e1c40a18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[138] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[139] = 80'h3f10a0b32f42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[139] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[140] = 80'hf8a042a8b1d1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[140] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[141] = 80'hc010041f98fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[141] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[142] = 80'h6f5155d6bf2a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[142] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[143] = 80'h6174e0aee88e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[143] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[144] = 80'hd8f296505931;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[144] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[145] = 80'he512e3c64789;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[145] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[146] = 80'h373e0b9976b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[146] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[147] = 80'h3e7dacda18b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[147] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[148] = 80'h964ddbc00a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[148] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[149] = 80'h54781b947c65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[149] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[150] = 80'h4e476ae23070;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[150] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[151] = 80'h965a202c5dd1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[151] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[152] = 80'h6eeef25e5a0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[152] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[153] = 80'hbd9be825e53c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[153] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[154] = 80'h5a0d2b0e2652;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[154] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[155] = 80'hf02c2960a78f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[155] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[156] = 80'h43801573ed5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[156] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[157] = 80'h34d1a3628645;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[157] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[158] = 80'h476d2c7ebc16;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[158] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[159] = 80'ha17de6c9b9c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[159] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[160] = 80'h2e3b2da7cb0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[160] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[161] = 80'h618fe75b3a00;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[161] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[162] = 80'h7868e9b929a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[162] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[163] = 80'hcbe5e4137d1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[163] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[164] = 80'h6771e8c490b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[164] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[165] = 80'h7be9cc15dbad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[165] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[166] = 80'h8c89b097b14c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[166] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[167] = 80'hf2124342ae18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[167] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[168] = 80'h330261ba3670;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[168] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[169] = 80'h42c4edb6d896;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[169] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[170] = 80'h23a570bc32da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[170] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[171] = 80'hdb4f2973fc73;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[171] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[172] = 80'h4c40d88318b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[172] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[173] = 80'h1273739101e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[173] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[174] = 80'h9c2ebac8770d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[174] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[175] = 80'haaeaffde1744;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[175] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[176] = 80'h67b1d0406ac4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[176] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[177] = 80'h602be7c25423;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[177] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[178] = 80'h7bd2374d89da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[178] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[179] = 80'h484efbf68ee5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[179] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[180] = 80'h8c2970d5df55;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[180] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[181] = 80'haec65cebfe7b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[181] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[182] = 80'h94dfc4cad63a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[182] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[183] = 80'h16398c9c5329;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[183] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[184] = 80'hc1d9c5b84501;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[184] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[185] = 80'hd1ad3332662b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[185] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[186] = 80'hb91d094ca5fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[186] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[187] = 80'h66807169ce5b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[187] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[188] = 80'h6ef096e4f564;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[188] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[189] = 80'h328864e675f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[189] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[190] = 80'h7dae2b0e1b45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[190] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[191] = 80'hbcb94b47b6e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[191] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[192] = 80'h969630df4be5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[192] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[193] = 80'h8fa1021a531a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[193] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[194] = 80'h872d61d5debf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[194] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[195] = 80'h991610788933;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[195] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[196] = 80'habf899e0a35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[196] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[197] = 80'h9a50b37b4c4e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[197] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[198] = 80'ha57859f9c477;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[198] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[199] = 80'h79cd60c49c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[199] = 80'h7fffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[200] = 80'h116a5a1abd7d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[200] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[201] = 80'hc21fd0b46818;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[201] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[202] = 80'hcb7c1d8cfffa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[202] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[203] = 80'h5da2668e789f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[203] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[204] = 80'ha975554d1660;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[204] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[205] = 80'hf527f8412a24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[205] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[206] = 80'h6e7cabe12a47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[206] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[207] = 80'hecce1c4cd86e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[207] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[208] = 80'h72d3d3fcd72b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[208] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[209] = 80'h839e1fb55d44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[209] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[210] = 80'h478398e0b9ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[210] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[211] = 80'h8530d50e759f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[211] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[212] = 80'h11f968361ebd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[212] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[213] = 80'h8ce994cc083f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[213] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[214] = 80'h2c23f84988ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[214] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[215] = 80'h9760938f25c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[215] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[216] = 80'h274efbfa8211;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[216] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[217] = 80'h694132b93ba3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[217] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[218] = 80'h682f3056401;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[218] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[219] = 80'hd1c36a785d4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[219] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[220] = 80'h4ae9b6d2ef4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[220] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[221] = 80'hc9c32ab41eeb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[221] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[222] = 80'hcbc076ebe28e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[222] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[223] = 80'hfbda31fd76c0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[223] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[224] = 80'h9a099a151b35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[224] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[225] = 80'h54a1681b3ffb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[225] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[226] = 80'hf0cf8f9ee272;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[226] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[227] = 80'h3f535b44d28a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[227] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[228] = 80'h7ae44fa333c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[228] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[229] = 80'hb665ce7f735a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[229] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[230] = 80'h626c7ae8774d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[230] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[231] = 80'hf3cddb51d392;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[231] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[232] = 80'h944a75a8319c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[232] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[233] = 80'heaacb9890fae;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[233] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[234] = 80'h46f6540ec7f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[234] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[235] = 80'hc6088fc1bd3d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[235] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[236] = 80'h5e0b61c56031;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[236] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[237] = 80'h27b4c51c3bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[237] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[238] = 80'hbe4d82d7e60e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[238] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[239] = 80'h7eef6a0932c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[239] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[240] = 80'h564f40cb3bc6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[240] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[241] = 80'h49ba0e14ede1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[241] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[242] = 80'hffa1385e8e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[242] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[243] = 80'hc2a6a6c5875c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[243] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[244] = 80'h46ed88992ff9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[244] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[245] = 80'h7bd52c488741;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[245] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[246] = 80'hdd037b320186;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[246] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[247] = 80'hbc45bae8ac0a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[247] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[248] = 80'h5b06c7e96f30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[248] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[249] = 80'hd4ddc557a673;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[249] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[250] = 80'h53ec21af6aa7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[250] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[251] = 80'h17ac57f88e87;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[251] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[252] = 80'ha4100e4032cc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[252] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[253] = 80'h140fa51dda60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[253] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[254] = 80'hba76b63b04af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[254] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[255] = 80'h7bf30212d42d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[255] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[256] = 80'h389a856d0929;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[256] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[257] = 80'h971def77bfa0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[257] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[258] = 80'h7fea6ca2dda9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[258] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[259] = 80'h6cc87b7163e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[259] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[260] = 80'h652f37432033;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[260] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[261] = 80'h94ca0afeaf40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[261] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[262] = 80'haa6075a82cfd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[262] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[263] = 80'he393132fbd4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[263] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[264] = 80'h8617fb8769a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[264] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[265] = 80'hd45704f554fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[265] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[266] = 80'h83aeac67707;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[266] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[267] = 80'had11dd592c9a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[267] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[268] = 80'h199fcd09ed28;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[268] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[269] = 80'h306fc67d4fd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[269] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[270] = 80'hded308236673;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[270] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[271] = 80'h6bb4f3981543;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[271] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[272] = 80'h28d774fa8bab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[272] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[273] = 80'h5f39e126fa40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[273] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[274] = 80'h4ec1930dd830;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[274] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[275] = 80'h2eabafa47444;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[275] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[276] = 80'hf2c4354979b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[276] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[277] = 80'h4375ff2839ff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[277] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[278] = 80'h831847d750e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[278] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[279] = 80'h6d4ff70a7fc3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[279] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[280] = 80'h67633ad96690;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[280] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[281] = 80'h58b1bb7ab35b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[281] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[282] = 80'h378d65b1297a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[282] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[283] = 80'h8ab24a720a34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[283] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[284] = 80'h9b617faf808a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[284] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[285] = 80'h2b5be33345f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[285] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[286] = 80'h80b069925240;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[286] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[287] = 80'h64819ae5ce38;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[287] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[288] = 80'hc8a2886319ad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[288] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[289] = 80'hbba80680cd74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[289] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[290] = 80'hc624c1780420;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[290] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[291] = 80'hdf4dc19f8a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[291] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[292] = 80'hbf4fc4c5109d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[292] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[293] = 80'h230e53a6e40d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[293] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[294] = 80'h6a8845704812;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[294] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[295] = 80'hd02d7e61c3ff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[295] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[296] = 80'h42d9ad4b7cb5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[296] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[297] = 80'h6620c43e40cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[297] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[298] = 80'h572b2a5075a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[298] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[299] = 80'hbc0a3cd8632;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[299] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[300] = 80'h318840f45c23;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[300] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[301] = 80'h7ec0b9f2df84;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[301] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[302] = 80'h708eaeea371;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[302] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[303] = 80'h29e3e9901c1f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[303] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[304] = 80'hf4f0fb40376f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[304] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[305] = 80'h7de8c27c7bf8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[305] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[306] = 80'h722214538bb3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[306] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[307] = 80'hb35284a2e8f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[307] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[308] = 80'hc1e963dc4088;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[308] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[309] = 80'h50d5503770e6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[309] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[310] = 80'hb63951662a30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[310] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[311] = 80'h7eddea567619;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[311] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[312] = 80'h4eab0a109e8f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[312] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[313] = 80'he549f26a551a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[313] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[314] = 80'h161e12d7d5f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[314] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[315] = 80'h2fb8691cf03d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[315] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[316] = 80'h6d0dd414bd88;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[316] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[317] = 80'hd47f0cfd8269;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[317] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[318] = 80'he7fe58f76aac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[318] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[319] = 80'hcddb5437e4b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[319] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[320] = 80'h58ac2d7d65c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[320] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[321] = 80'he81d8eb85034;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[321] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[322] = 80'ha6fb99d69d1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[322] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[323] = 80'h85db0f2ad52e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[323] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[324] = 80'hba447f49c0b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[324] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[325] = 80'h99d3496acd35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[325] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[326] = 80'h40e7e1b07303;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[326] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[327] = 80'h55f948ebe91d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[327] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[328] = 80'h392c0459ce02;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[328] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[329] = 80'h7e3d419f5d34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[329] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[330] = 80'he74efb58eaa7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[330] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[331] = 80'hf83f581e4482;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[331] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[332] = 80'h9cce1dfeef14;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[332] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[333] = 80'h4b70936e9f64;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[333] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[334] = 80'h8f60bf446783;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[334] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[335] = 80'h93a9046448e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[335] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[336] = 80'h6e3ce4ac6730;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[336] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[337] = 80'h84de22fbc40a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[337] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[338] = 80'h2d98732c0914;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[338] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[339] = 80'h588e0584287c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[339] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[340] = 80'h8f50e0497e89;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[340] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[341] = 80'hb0e119fb2555;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[341] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[342] = 80'h4cd3c2cde21a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[342] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[343] = 80'hda342cb3beee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[343] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[344] = 80'h9f7fc5e6a042;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[344] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[345] = 80'hcc5300c82669;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[345] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[346] = 80'h6a1ec386bf00;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[346] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[347] = 80'h2317e8d90545;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[347] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[348] = 80'h8d4fe98625cf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[348] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[349] = 80'h60665e2c19e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[349] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[350] = 80'h596674fbbfb1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[350] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[351] = 80'h5c7688d8aad5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[351] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[352] = 80'h99c3cb202d30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[352] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[353] = 80'ha86ac83a7681;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[353] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[354] = 80'hf9f330aaf7e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[354] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[355] = 80'h3c3dcdb988e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[355] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[356] = 80'h82440e73e0a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[356] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[357] = 80'hdeb63d376bdd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[357] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[358] = 80'h3f13c6d986da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[358] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[359] = 80'h959a11161a8a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[359] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[360] = 80'h4fc4b9709a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[360] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[361] = 80'h603260a4fa8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[361] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[362] = 80'h317642426d30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[362] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[363] = 80'h93eea5159da0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[363] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[364] = 80'ha6a6c5effbb8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[364] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[365] = 80'h9a556fc0f1e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[365] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[366] = 80'hca8bfde422b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[366] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[367] = 80'h6b3d4da4a0e4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[367] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[368] = 80'hb8725432eee0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[368] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[369] = 80'h2a5f4d97572c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[369] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[370] = 80'h3f4b2f37c91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[370] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[371] = 80'h6d012a56f306;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[371] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[372] = 80'hf39c18ff7423;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[372] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[373] = 80'h64fe54c3d020;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[373] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[374] = 80'h5941386df853;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[374] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[375] = 80'hfd5081a7023d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[375] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[376] = 80'h59d252677e44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[376] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[377] = 80'hb1ef710456c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[377] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[378] = 80'h8a3b29afa55f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[378] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[379] = 80'ha8f4af7c920a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[379] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[380] = 80'h9b5b556528f0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[380] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[381] = 80'h8d75c4ce6384;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[381] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[382] = 80'h644e172a4d39;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[382] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[383] = 80'h4e2c31c4e9bf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[383] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[384] = 80'hfb16e104670e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[384] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[385] = 80'hedda66338267;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[385] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[386] = 80'h28c12a16f1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[386] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[387] = 80'hff84824ad314;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[387] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[388] = 80'hbe7756aeeab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[388] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[389] = 80'h7e61e055303f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[389] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[390] = 80'haac7193a22af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[390] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[391] = 80'h565f0106873e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[391] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[392] = 80'h75032e61802d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[392] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[393] = 80'hf2f7c9dbbf6e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[393] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[394] = 80'hc616b82074dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[394] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[395] = 80'h9b90c73a26b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[395] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[396] = 80'hf1aad48501e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[396] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[397] = 80'hb50e5a5b2331;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[397] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[398] = 80'h536e70ff511;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[398] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[399] = 80'h500f137223d6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[399] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[400] = 80'h2791051b62a6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[400] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[401] = 80'hc4eb2c045df0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[401] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[402] = 80'ha4ad1b4e4c65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[402] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[403] = 80'h5dcd203c62ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[403] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[404] = 80'hbd2053fe1aa1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[404] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[405] = 80'hdd873733eebd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[405] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[406] = 80'hd5cc8944cc44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[406] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[407] = 80'hdf75e34c1d60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[407] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[408] = 80'h69516c90e02b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[408] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[409] = 80'hba7434218648;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[409] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[410] = 80'h75995e082cc9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[410] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[411] = 80'h8f8a0618c492;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[411] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[412] = 80'h85652adefb50;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[412] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[413] = 80'h84e3bbb346a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[413] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[414] = 80'hce288545ff5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[414] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[415] = 80'hf34840529bc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[415] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[416] = 80'h93b680734ca8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[416] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[417] = 80'h6d3e5930bf31;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[417] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[418] = 80'h4c6bb4e13dd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[418] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[419] = 80'hc17e7cae146d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[419] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[420] = 80'h3a01e234f448;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[420] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[421] = 80'h1f6089a70d31;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[421] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[422] = 80'he9910acedf01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[422] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[423] = 80'h92c1be63a45c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[423] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[424] = 80'h77250b5545e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[424] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[425] = 80'h41875a4af1b4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[425] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[426] = 80'h1f7188b8f195;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[426] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[427] = 80'he7043697f5e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[427] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[428] = 80'hccb0a5325cbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[428] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[429] = 80'hf77c99d0ae10;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[429] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[430] = 80'h51c66267cec7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[430] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[431] = 80'ha3eb7b517f7d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[431] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[432] = 80'h5e4b84a9a324;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[432] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[433] = 80'h263366d9a934;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[433] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[434] = 80'h35cd167e2bad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[434] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[435] = 80'hb2c3bbf8fba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[435] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[436] = 80'h8f19a66976c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[436] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[437] = 80'he0b42c35622b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[437] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[438] = 80'hdca9a6f1782c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[438] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[439] = 80'h9a1541c274a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[439] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[440] = 80'h44768a38b95d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[440] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[441] = 80'h38f48a68b142;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[441] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[442] = 80'h9759c188b4fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[442] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[443] = 80'ha08c0f3399b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[443] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[444] = 80'h820dea118ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[444] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[445] = 80'h786f4fec3569;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[445] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[446] = 80'h35502a9bf339;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[446] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[447] = 80'hede032f81911;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[447] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[448] = 80'h5d2da41d57;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[448] = 80'h7fffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[449] = 80'h1d551e45233a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[449] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[450] = 80'h1232e7e21619;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[450] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[451] = 80'h9656bf8e0b9d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[451] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[452] = 80'h282df63c9a42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[452] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[453] = 80'hfb8cfa3efc1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[453] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[454] = 80'he202a5e04142;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[454] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[455] = 80'hce14bd93ed55;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[455] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[456] = 80'hb29b6b75332;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[456] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[457] = 80'ha560cfe7acfc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[457] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[458] = 80'h99c7f0448e01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[458] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[459] = 80'h1dc007e9c85a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[459] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[460] = 80'hd5bbfcebded1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[460] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[461] = 80'h7a59ce859cc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[461] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[462] = 80'h4ea8c5b70bda;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[462] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[463] = 80'h52f1807fc08a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[463] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[464] = 80'h206171d9529a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[464] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[465] = 80'h498a7ea9d6a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[465] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[466] = 80'h68b1d8990008;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[466] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[467] = 80'hdfdd7f5c6649;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[467] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[468] = 80'h423c83f43d47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[468] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[469] = 80'h71daa74440c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[469] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[470] = 80'h6b7caeb2cb69;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[470] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[471] = 80'h9301716b199f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[471] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[472] = 80'hf30c2c261355;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[472] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[473] = 80'he1037b5789b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[473] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[474] = 80'h4ac85c163c30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[474] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[475] = 80'hbd2e17a3bd71;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[475] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[476] = 80'h8cfbaac12a25;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[476] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[477] = 80'he07f86b355a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[477] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[478] = 80'he24b3b5f435d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[478] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[479] = 80'hc6100a3221e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[479] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[480] = 80'hd601e9e5d6ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[480] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[481] = 80'ha2ee82f9007b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[481] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[482] = 80'hb4baf8944204;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[482] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[483] = 80'h78c5ee1f506d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[483] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[484] = 80'h94176a64d950;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[484] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[485] = 80'hbdc7edf2bed3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[485] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[486] = 80'hf6141087125a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[486] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[487] = 80'h4d8a6c4bb175;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[487] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[488] = 80'hd702b7ff755e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[488] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[489] = 80'h17ad459c4491;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[489] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[490] = 80'hbecd69de0af5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[490] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[491] = 80'h6db83a09cb40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[491] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[492] = 80'hc15a3192c54e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[492] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[493] = 80'h372729de79a7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[493] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[494] = 80'hb7d5a573112e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[494] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[495] = 80'he7598a8d64ef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[495] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[496] = 80'h4d77a8f186e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[496] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[497] = 80'hb3a7e8c62438;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[497] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[498] = 80'h5e628e40bad8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[498] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[499] = 80'h2c6ae9566a81;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[499] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[500] = 80'h7c8088a4d780;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[500] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[501] = 80'h449da718991b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[501] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[502] = 80'heb14915c851e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[502] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[503] = 80'h3527b3d245b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[503] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[504] = 80'h85d7cc131a8a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[504] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[505] = 80'hb448dcc734b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[505] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[506] = 80'h463282aaf56;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[506] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[507] = 80'he6f6fe35b667;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[507] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[508] = 80'h80c258b15826;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[508] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[509] = 80'hfaac4f7283f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[509] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[510] = 80'ha03cce697a88;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[510] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[511] = 80'hdf03c7e186d0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[511] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[512] = 80'hc301b2ddb491;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[512] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[513] = 80'h5a553a6d946;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[513] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[514] = 80'hec81a0ecf565;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[514] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[515] = 80'h25b7ba6c7a22;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[515] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[516] = 80'hff62f77af68e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[516] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[517] = 80'h90696c0e7c49;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[517] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[518] = 80'hdb542752b51b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[518] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[519] = 80'h5c669d7e5719;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[519] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[520] = 80'h7869b90d6d6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[520] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[521] = 80'h6ab3f4028bc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[521] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[522] = 80'hfaf254c81784;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[522] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[523] = 80'he91e80ddf2b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[523] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[524] = 80'h12ec8002dccf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[524] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[525] = 80'h1fb66119b301;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[525] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[526] = 80'h35cfa56dca6a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[526] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[527] = 80'h257f17287640;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[527] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[528] = 80'he24b719e5fd5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[528] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[529] = 80'h1b6de98d63bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[529] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[530] = 80'hc7396a1e1d0b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[530] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[531] = 80'h7fb43ae9cd4b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[531] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[532] = 80'ha389a8825008;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[532] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[533] = 80'h62002cc089d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[533] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[534] = 80'ha2fc3e097fd8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[534] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[535] = 80'h93938f2e7bb6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[535] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[536] = 80'h4c0878c8f3c9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[536] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[537] = 80'h6dad4681d74b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[537] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[538] = 80'h90d849afd440;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[538] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[539] = 80'h99cea5c192b2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[539] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[540] = 80'h439a63924ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[540] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[541] = 80'h22efe4c3db4e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[541] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[542] = 80'h935f8ae1eaca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[542] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[543] = 80'h980ce89cb3ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[543] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[544] = 80'hb2b1d54e6143;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[544] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[545] = 80'h985262ca09c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[545] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[546] = 80'h1b5370c23148;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[546] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[547] = 80'hfa6e44897737;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[547] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[548] = 80'hedc347b5f551;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[548] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[549] = 80'hbbafbcb86844;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[549] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[550] = 80'h7fb9ba95cb59;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[550] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[551] = 80'hbe931b35ee21;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[551] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[552] = 80'h39f56d709e34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[552] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[553] = 80'h4e9dfa08200a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[553] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[554] = 80'h820c31b21a45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[554] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[555] = 80'h5c7809f7005;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[555] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[556] = 80'h3aca0c094cca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[556] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[557] = 80'h745ae42f60b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[557] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[558] = 80'h9ab1034e7c6e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[558] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[559] = 80'h8b03e00b02c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[559] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[560] = 80'h291393c268aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[560] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[561] = 80'h4f5dda910b46;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[561] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[562] = 80'hd702572b740;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[562] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[563] = 80'h82eb751a50eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[563] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[564] = 80'h69f1bf212be5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[564] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[565] = 80'h692f8eeae2e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[565] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[566] = 80'h19a683169415;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[566] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[567] = 80'h93bac3e6e685;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[567] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[568] = 80'h4993bee769ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[568] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[569] = 80'hcd7fb4cb6753;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[569] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[570] = 80'h240e7a3c36d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[570] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[571] = 80'hdee7cb29be85;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[571] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[572] = 80'h992597565e42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[572] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[573] = 80'h5cf48819c736;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[573] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[574] = 80'h47abe210da7f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[574] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[575] = 80'hf93a1757baa0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[575] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[576] = 80'h7c1ceb4afc56;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[576] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[577] = 80'haf7d256d7cc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[577] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[578] = 80'h56f4eacb32c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[578] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[579] = 80'hb0d1add53e47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[579] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[580] = 80'hd2755cc4bd17;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[580] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[581] = 80'ha6985589f9f2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[581] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[582] = 80'hc617a79d7ece;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[582] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[583] = 80'hce74602fffba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[583] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[584] = 80'hf924b4b96d61;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[584] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[585] = 80'h8c0b6b9901dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[585] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[586] = 80'hf68af87708bf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[586] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[587] = 80'h74fa5f30fe3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[587] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[588] = 80'h4db8a921b1d2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[588] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[589] = 80'h18a72f979e24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[589] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[590] = 80'h595e18260e26;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[590] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[591] = 80'haad2d483e822;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[591] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[592] = 80'h343913fad305;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[592] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[593] = 80'hb3d2b6c10e97;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[593] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[594] = 80'h5b359f4f70b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[594] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[595] = 80'h910fdf65238e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[595] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[596] = 80'h858d2a03d342;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[596] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[597] = 80'h60c0b6079327;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[597] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[598] = 80'hac7bf03559d7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[598] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[599] = 80'h9ad2390bbe32;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[599] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[600] = 80'hfa4f7ce06718;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[600] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[601] = 80'hd16fe65ec39f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[601] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[602] = 80'h2d99e55053a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[602] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[603] = 80'h5159029f3697;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[603] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[604] = 80'hb4b0447b5549;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[604] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[605] = 80'h377b752a37b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[605] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[606] = 80'h220bb11437f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[606] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[607] = 80'habd69fb1204e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[607] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[608] = 80'heb47988d0d8b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[608] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[609] = 80'hca9cc767edce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[609] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[610] = 80'h3b6f42cbe0a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[610] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[611] = 80'h1dd3fa287076;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[611] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[612] = 80'h9628912dbff2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[612] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[613] = 80'h89a7951bea35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[613] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[614] = 80'hc7b2ff90ab75;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[614] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[615] = 80'h7ec37d3f35d1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[615] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[616] = 80'h486d45350ba4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[616] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[617] = 80'hf7c78a4aeffd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[617] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[618] = 80'hea7f3c4470a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[618] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[619] = 80'h95398bca46db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[619] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[620] = 80'h2a21d269ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[620] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[621] = 80'h5ff142432afa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[621] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[622] = 80'h8d346fc65e2b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[622] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[623] = 80'h1a6584f50556;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[623] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[624] = 80'h8386da1029f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[624] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[625] = 80'hdb56c981ece6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[625] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[626] = 80'hcfe8af38f522;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[626] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[627] = 80'h8e919d8a745b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[627] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[628] = 80'h543818958c78;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[628] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[629] = 80'ha8b931f97188;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[629] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[630] = 80'h7dee0d849922;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[630] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[631] = 80'h1017ca8a2953;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[631] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[632] = 80'h7ed9cae24403;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[632] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[633] = 80'hea187ed4d55a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[633] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[634] = 80'h2e76e28270f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[634] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[635] = 80'hf1980343333f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[635] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[636] = 80'h8de1c963c062;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[636] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[637] = 80'h3fd86ea44501;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[637] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[638] = 80'hdc791a00bf2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[638] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[639] = 80'h76fd772b3105;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[639] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[640] = 80'h9137a6d429b2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[640] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[641] = 80'h49d4cbef7ccc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[641] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[642] = 80'h8051f12b529f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[642] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[643] = 80'h8d6aa657a5e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[643] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[644] = 80'h44bafb829ee6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[644] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[645] = 80'he55061ccc7b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[645] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[646] = 80'hd75970bd3bb0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[646] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[647] = 80'h4811729ba385;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[647] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[648] = 80'hc0501fd955df;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[648] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[649] = 80'h659c29b06d69;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[649] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[650] = 80'h6aec373261a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[650] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[651] = 80'hc25cd90f5dab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[651] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[652] = 80'hcee3230bfef6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[652] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[653] = 80'h7bde198a992f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[653] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[654] = 80'h7cd4d9587ccb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[654] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[655] = 80'h5cee7e94dd42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[655] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[656] = 80'hc7f2c96b613;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[656] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[657] = 80'hf2de9d0bdde4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[657] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[658] = 80'hb80342294761;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[658] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[659] = 80'hef05f9051dde;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[659] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[660] = 80'h89d9864b0f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[660] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[661] = 80'hf84ebc6b5933;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[661] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[662] = 80'h99c7ebd6ef11;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[662] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[663] = 80'ha5cfc726453c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[663] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[664] = 80'h8e33ccc43905;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[664] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[665] = 80'h61dbc393f8b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[665] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[666] = 80'hb5776eb8e40c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[666] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[667] = 80'hc56f02fbb8af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[667] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[668] = 80'hf06ac89a6e2e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[668] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[669] = 80'h4d46ea5704c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[669] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[670] = 80'h18a0d2ab536;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[670] = 80'h1ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[671] = 80'hde24ea9c8559;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[671] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[672] = 80'h117c2dcb8a3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[672] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[673] = 80'h42c5800a198;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[673] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[674] = 80'hc866641162c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[674] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[675] = 80'hc59ce2a178ef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[675] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[676] = 80'h91b9a88b2186;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[676] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[677] = 80'hbaaaa92f9330;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[677] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[678] = 80'h899bc4d45fed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[678] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[679] = 80'h31aba86c07cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[679] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[680] = 80'hc4984e56b9a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[680] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[681] = 80'h1b2cb5378bd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[681] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[682] = 80'hff120ca68f9a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[682] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[683] = 80'ha835dfd4a64e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[683] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[684] = 80'hcc35683c57dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[684] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[685] = 80'ha5c1099a0ccc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[685] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[686] = 80'hefd95c4e5fe9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[686] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[687] = 80'h7c76d25796aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[687] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[688] = 80'h7b60730923d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[688] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[689] = 80'h7373b8b8f3c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[689] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[690] = 80'h37e56c799b77;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[690] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[691] = 80'h64aeec7ab84c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[691] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[692] = 80'hdc1814387312;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[692] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[693] = 80'hdd2835b8c4f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[693] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[694] = 80'h5af2eb552cca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[694] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[695] = 80'h446b9299fa74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[695] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[696] = 80'h86928cf64fc6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[696] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[697] = 80'hc4fdc019c61f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[697] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[698] = 80'h882f97bb161f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[698] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[699] = 80'h4ed606f4518d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[699] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem[700] = 80'hbd46a3aa3c15;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[2].u_tcam.mem_mask[700] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[0] = 80'h0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[1] = 80'hc76428a3ac18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[1] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[2] = 80'h6fa2b332a044;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[2] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[3] = 80'hdf160ea7e244;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[3] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[4] = 80'hbde8a5158a2b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[4] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[5] = 80'h1c7fcaa5772f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[5] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[6] = 80'h398bc2065413;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[6] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[7] = 80'hbf26a132d23e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[7] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[8] = 80'h2e5a52ddfb3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[8] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[9] = 80'hf9c4f448c4c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[9] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[10] = 80'h35e4dd182f90;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[10] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[11] = 80'h8513d0c50521;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[11] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[12] = 80'h35a66285b62e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[12] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[13] = 80'h4915d9de428f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[13] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[14] = 80'h3eff489073c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[14] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[15] = 80'hd00165db49c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[15] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[16] = 80'hc6e7d540048a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[16] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[17] = 80'hd2cf31221e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[17] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[18] = 80'h9cc2400c08bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[18] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[19] = 80'he84ab68b1a24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[19] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[20] = 80'hdc9c606e91ae;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[20] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[21] = 80'h4b8ee53f7660;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[21] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[22] = 80'ha6dc109cdbbd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[22] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[23] = 80'h2e5acd726cb2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[23] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[24] = 80'hbb30b2ecd487;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[24] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[25] = 80'h9aeec82f8fac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[25] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[26] = 80'hab83fe2b985c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[26] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[27] = 80'hca3daac02b2f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[27] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[28] = 80'h1a893b2ffa10;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[28] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[29] = 80'hcb1ab883d9ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[29] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[30] = 80'h6ddb0412e88d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[30] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[31] = 80'h25d034a677c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[31] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[32] = 80'h2ee63ce89af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[32] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[33] = 80'h1ab5a710d843;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[33] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[34] = 80'h97e8c062f084;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[34] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[35] = 80'h30a809743d4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[35] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[36] = 80'h22420da7f8f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[36] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[37] = 80'hafaf284ad3bc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[37] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[38] = 80'h53bd4f0d7794;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[38] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[39] = 80'h5c0d39f2f061;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[39] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[40] = 80'h9419a7ce074a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[40] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[41] = 80'h52d45cc1e4a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[41] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[42] = 80'h9b30665b9971;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[42] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[43] = 80'h20d936f412c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[43] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[44] = 80'h8b889af41550;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[44] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[45] = 80'hf91ce85e797d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[45] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[46] = 80'h6e1dbd81191;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[46] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[47] = 80'h345e3c5f1365;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[47] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[48] = 80'h8dceefe91dc9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[48] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[49] = 80'hd47d2191ffed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[49] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[50] = 80'h7d341fbc821b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[50] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[51] = 80'h2e1c5d9ff7d9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[51] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[52] = 80'hb7c667fd0324;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[52] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[53] = 80'h4933bf21a16c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[53] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[54] = 80'hf9724902347e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[54] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[55] = 80'haeb766b220db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[55] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[56] = 80'hdbbc2a3224ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[56] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[57] = 80'h365a679e8085;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[57] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[58] = 80'heeff7c2b7b33;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[58] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[59] = 80'h45bb6a31bb68;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[59] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[60] = 80'h1a81b1c43f91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[60] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[61] = 80'h1de0ad29184a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[61] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[62] = 80'h4eb9229cd415;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[62] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[63] = 80'h75c39cfd15db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[63] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[64] = 80'hbd7d9ddf726;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[64] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[65] = 80'h788ece7eed43;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[65] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[66] = 80'h689790000fff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[66] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[67] = 80'h30fca31cf96b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[67] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[68] = 80'h358975cc2823;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[68] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[69] = 80'h6b1cd921c79d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[69] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[70] = 80'h549a31ff63b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[70] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[71] = 80'h310dee607220;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[71] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[72] = 80'haf90fc2fb606;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[72] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[73] = 80'hdb655000d3a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[73] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[74] = 80'h8bf35344ab45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[74] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[75] = 80'h2d8a38190b20;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[75] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[76] = 80'h263f7f66582;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[76] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[77] = 80'h4dfc2ba4768d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[77] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[78] = 80'h849983bfbe7a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[78] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[79] = 80'h1efcb2f4dd4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[79] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[80] = 80'h61e5a9de4569;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[80] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[81] = 80'h770c1c4bd3a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[81] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[82] = 80'h500562660aff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[82] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[83] = 80'ha72a189143e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[83] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[84] = 80'h51a64abf0e09;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[84] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[85] = 80'h1f5700abe928;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[85] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[86] = 80'h512e72fad6a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[86] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[87] = 80'h5f3a530396cf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[87] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[88] = 80'h748487400445;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[88] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[89] = 80'h87719fb3f864;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[89] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[90] = 80'he88c8f60061d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[90] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[91] = 80'h9f6cc5f93019;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[91] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[92] = 80'hfa9df2c0fa11;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[92] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[93] = 80'h3e5de237f4f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[93] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[94] = 80'h1220e6f8b9fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[94] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[95] = 80'hceb0c2f94c3c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[95] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[96] = 80'h1845b8356ded;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[96] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[97] = 80'hcb7d6f052ed9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[97] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[98] = 80'ha1d827523dc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[98] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[99] = 80'hcaf8264a3ea;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[99] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[100] = 80'h38ead3f12916;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[100] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[101] = 80'h13d2ee37c448;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[101] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[102] = 80'h3c2fe7d9f34c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[102] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[103] = 80'h3c1db8626079;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[103] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[104] = 80'h865b861ca607;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[104] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[105] = 80'h794600c6d0f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[105] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[106] = 80'he00c57f6e0b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[106] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[107] = 80'he29db65e8903;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[107] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[108] = 80'h8e261e6170f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[108] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[109] = 80'h66939b10ec73;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[109] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[110] = 80'h70c2e9c3c8eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[110] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[111] = 80'h45c66be84cf4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[111] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[112] = 80'h232cef211d0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[112] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[113] = 80'h80542dda5aa2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[113] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[114] = 80'h474effbc30dd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[114] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[115] = 80'he4cebd5c6fa4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[115] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[116] = 80'haf6a54830375;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[116] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[117] = 80'h8ef028be44c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[117] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[118] = 80'h5fdca8436bf4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[118] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[119] = 80'h6e7e1c15bd08;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[119] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[120] = 80'h134c1f65fd66;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[120] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[121] = 80'hcea87493679f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[121] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[122] = 80'hceb7bc309c1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[122] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[123] = 80'h61a6f8771878;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[123] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[124] = 80'hcedef6a567fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[124] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[125] = 80'h2e32a08622cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[125] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[126] = 80'h5356e16b8fd7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[126] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[127] = 80'hfd605bd942c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[127] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[128] = 80'hd5f103f449;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[128] = 80'hffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[129] = 80'h5f57f4362b22;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[129] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[130] = 80'h2e67f284f871;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[130] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[131] = 80'hecd79dcadc01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[131] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[132] = 80'he00525c7b0f8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[132] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[133] = 80'hb3cf483e6c80;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[133] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[134] = 80'h77eb26f31bbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[134] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[135] = 80'h8b676c49d915;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[135] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[136] = 80'ha2822acbd35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[136] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[137] = 80'h3a257929df1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[137] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[138] = 80'he9b0e1c40a18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[138] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[139] = 80'h3f10a0b32f42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[139] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[140] = 80'hf8a042a8b1d1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[140] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[141] = 80'hc010041f98fe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[141] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[142] = 80'h6f5155d6bf2a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[142] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[143] = 80'h6174e0aee88e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[143] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[144] = 80'hd8f296505931;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[144] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[145] = 80'he512e3c64789;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[145] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[146] = 80'h373e0b9976b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[146] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[147] = 80'h3e7dacda18b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[147] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[148] = 80'h964ddbc00a5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[148] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[149] = 80'h54781b947c65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[149] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[150] = 80'h4e476ae23070;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[150] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[151] = 80'h965a202c5dd1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[151] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[152] = 80'h6eeef25e5a0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[152] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[153] = 80'hbd9be825e53c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[153] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[154] = 80'h5a0d2b0e2652;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[154] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[155] = 80'hf02c2960a78f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[155] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[156] = 80'h43801573ed5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[156] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[157] = 80'h34d1a3628645;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[157] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[158] = 80'h476d2c7ebc16;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[158] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[159] = 80'ha17de6c9b9c6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[159] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[160] = 80'h2e3b2da7cb0e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[160] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[161] = 80'h618fe75b3a00;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[161] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[162] = 80'h7868e9b929a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[162] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[163] = 80'hcbe5e4137d1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[163] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[164] = 80'h6771e8c490b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[164] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[165] = 80'h7be9cc15dbad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[165] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[166] = 80'h8c89b097b14c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[166] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[167] = 80'hf2124342ae18;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[167] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[168] = 80'h330261ba3670;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[168] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[169] = 80'h42c4edb6d896;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[169] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[170] = 80'h23a570bc32da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[170] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[171] = 80'hdb4f2973fc73;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[171] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[172] = 80'h4c40d88318b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[172] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[173] = 80'h1273739101e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[173] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[174] = 80'h9c2ebac8770d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[174] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[175] = 80'haaeaffde1744;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[175] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[176] = 80'h67b1d0406ac4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[176] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[177] = 80'h602be7c25423;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[177] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[178] = 80'h7bd2374d89da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[178] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[179] = 80'h484efbf68ee5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[179] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[180] = 80'h8c2970d5df55;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[180] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[181] = 80'haec65cebfe7b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[181] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[182] = 80'h94dfc4cad63a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[182] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[183] = 80'h16398c9c5329;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[183] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[184] = 80'hc1d9c5b84501;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[184] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[185] = 80'hd1ad3332662b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[185] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[186] = 80'hb91d094ca5fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[186] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[187] = 80'h66807169ce5b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[187] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[188] = 80'h6ef096e4f564;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[188] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[189] = 80'h328864e675f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[189] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[190] = 80'h7dae2b0e1b45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[190] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[191] = 80'hbcb94b47b6e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[191] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[192] = 80'h969630df4be5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[192] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[193] = 80'h8fa1021a531a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[193] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[194] = 80'h872d61d5debf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[194] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[195] = 80'h991610788933;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[195] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[196] = 80'habf899e0a35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[196] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[197] = 80'h9a50b37b4c4e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[197] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[198] = 80'ha57859f9c477;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[198] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[199] = 80'h79cd60c49c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[199] = 80'h7fffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[200] = 80'h116a5a1abd7d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[200] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[201] = 80'hc21fd0b46818;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[201] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[202] = 80'hcb7c1d8cfffa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[202] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[203] = 80'h5da2668e789f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[203] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[204] = 80'ha975554d1660;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[204] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[205] = 80'hf527f8412a24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[205] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[206] = 80'h6e7cabe12a47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[206] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[207] = 80'hecce1c4cd86e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[207] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[208] = 80'h72d3d3fcd72b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[208] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[209] = 80'h839e1fb55d44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[209] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[210] = 80'h478398e0b9ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[210] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[211] = 80'h8530d50e759f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[211] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[212] = 80'h11f968361ebd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[212] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[213] = 80'h8ce994cc083f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[213] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[214] = 80'h2c23f84988ee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[214] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[215] = 80'h9760938f25c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[215] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[216] = 80'h274efbfa8211;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[216] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[217] = 80'h694132b93ba3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[217] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[218] = 80'h682f3056401;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[218] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[219] = 80'hd1c36a785d4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[219] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[220] = 80'h4ae9b6d2ef4f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[220] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[221] = 80'hc9c32ab41eeb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[221] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[222] = 80'hcbc076ebe28e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[222] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[223] = 80'hfbda31fd76c0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[223] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[224] = 80'h9a099a151b35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[224] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[225] = 80'h54a1681b3ffb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[225] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[226] = 80'hf0cf8f9ee272;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[226] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[227] = 80'h3f535b44d28a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[227] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[228] = 80'h7ae44fa333c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[228] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[229] = 80'hb665ce7f735a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[229] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[230] = 80'h626c7ae8774d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[230] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[231] = 80'hf3cddb51d392;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[231] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[232] = 80'h944a75a8319c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[232] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[233] = 80'heaacb9890fae;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[233] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[234] = 80'h46f6540ec7f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[234] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[235] = 80'hc6088fc1bd3d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[235] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[236] = 80'h5e0b61c56031;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[236] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[237] = 80'h27b4c51c3bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[237] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[238] = 80'hbe4d82d7e60e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[238] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[239] = 80'h7eef6a0932c5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[239] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[240] = 80'h564f40cb3bc6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[240] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[241] = 80'h49ba0e14ede1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[241] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[242] = 80'hffa1385e8e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[242] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[243] = 80'hc2a6a6c5875c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[243] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[244] = 80'h46ed88992ff9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[244] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[245] = 80'h7bd52c488741;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[245] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[246] = 80'hdd037b320186;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[246] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[247] = 80'hbc45bae8ac0a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[247] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[248] = 80'h5b06c7e96f30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[248] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[249] = 80'hd4ddc557a673;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[249] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[250] = 80'h53ec21af6aa7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[250] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[251] = 80'h17ac57f88e87;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[251] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[252] = 80'ha4100e4032cc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[252] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[253] = 80'h140fa51dda60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[253] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[254] = 80'hba76b63b04af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[254] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[255] = 80'h7bf30212d42d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[255] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[256] = 80'h389a856d0929;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[256] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[257] = 80'h971def77bfa0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[257] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[258] = 80'h7fea6ca2dda9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[258] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[259] = 80'h6cc87b7163e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[259] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[260] = 80'h652f37432033;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[260] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[261] = 80'h94ca0afeaf40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[261] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[262] = 80'haa6075a82cfd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[262] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[263] = 80'he393132fbd4d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[263] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[264] = 80'h8617fb8769a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[264] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[265] = 80'hd45704f554fa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[265] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[266] = 80'h83aeac67707;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[266] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[267] = 80'had11dd592c9a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[267] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[268] = 80'h199fcd09ed28;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[268] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[269] = 80'h306fc67d4fd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[269] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[270] = 80'hded308236673;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[270] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[271] = 80'h6bb4f3981543;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[271] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[272] = 80'h28d774fa8bab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[272] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[273] = 80'h5f39e126fa40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[273] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[274] = 80'h4ec1930dd830;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[274] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[275] = 80'h2eabafa47444;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[275] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[276] = 80'hf2c4354979b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[276] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[277] = 80'h4375ff2839ff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[277] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[278] = 80'h831847d750e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[278] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[279] = 80'h6d4ff70a7fc3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[279] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[280] = 80'h67633ad96690;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[280] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[281] = 80'h58b1bb7ab35b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[281] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[282] = 80'h378d65b1297a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[282] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[283] = 80'h8ab24a720a34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[283] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[284] = 80'h9b617faf808a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[284] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[285] = 80'h2b5be33345f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[285] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[286] = 80'h80b069925240;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[286] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[287] = 80'h64819ae5ce38;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[287] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[288] = 80'hc8a2886319ad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[288] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[289] = 80'hbba80680cd74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[289] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[290] = 80'hc624c1780420;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[290] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[291] = 80'hdf4dc19f8a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[291] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[292] = 80'hbf4fc4c5109d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[292] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[293] = 80'h230e53a6e40d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[293] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[294] = 80'h6a8845704812;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[294] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[295] = 80'hd02d7e61c3ff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[295] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[296] = 80'h42d9ad4b7cb5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[296] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[297] = 80'h6620c43e40cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[297] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[298] = 80'h572b2a5075a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[298] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[299] = 80'hbc0a3cd8632;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[299] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[300] = 80'h318840f45c23;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[300] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[301] = 80'h7ec0b9f2df84;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[301] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[302] = 80'h708eaeea371;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[302] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[303] = 80'h29e3e9901c1f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[303] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[304] = 80'hf4f0fb40376f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[304] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[305] = 80'h7de8c27c7bf8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[305] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[306] = 80'h722214538bb3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[306] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[307] = 80'hb35284a2e8f3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[307] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[308] = 80'hc1e963dc4088;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[308] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[309] = 80'h50d5503770e6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[309] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[310] = 80'hb63951662a30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[310] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[311] = 80'h7eddea567619;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[311] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[312] = 80'h4eab0a109e8f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[312] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[313] = 80'he549f26a551a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[313] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[314] = 80'h161e12d7d5f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[314] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[315] = 80'h2fb8691cf03d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[315] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[316] = 80'h6d0dd414bd88;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[316] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[317] = 80'hd47f0cfd8269;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[317] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[318] = 80'he7fe58f76aac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[318] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[319] = 80'hcddb5437e4b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[319] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[320] = 80'h58ac2d7d65c1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[320] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[321] = 80'he81d8eb85034;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[321] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[322] = 80'ha6fb99d69d1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[322] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[323] = 80'h85db0f2ad52e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[323] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[324] = 80'hba447f49c0b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[324] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[325] = 80'h99d3496acd35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[325] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[326] = 80'h40e7e1b07303;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[326] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[327] = 80'h55f948ebe91d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[327] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[328] = 80'h392c0459ce02;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[328] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[329] = 80'h7e3d419f5d34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[329] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[330] = 80'he74efb58eaa7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[330] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[331] = 80'hf83f581e4482;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[331] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[332] = 80'h9cce1dfeef14;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[332] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[333] = 80'h4b70936e9f64;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[333] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[334] = 80'h8f60bf446783;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[334] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[335] = 80'h93a9046448e2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[335] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[336] = 80'h6e3ce4ac6730;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[336] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[337] = 80'h84de22fbc40a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[337] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[338] = 80'h2d98732c0914;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[338] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[339] = 80'h588e0584287c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[339] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[340] = 80'h8f50e0497e89;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[340] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[341] = 80'hb0e119fb2555;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[341] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[342] = 80'h4cd3c2cde21a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[342] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[343] = 80'hda342cb3beee;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[343] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[344] = 80'h9f7fc5e6a042;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[344] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[345] = 80'hcc5300c82669;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[345] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[346] = 80'h6a1ec386bf00;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[346] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[347] = 80'h2317e8d90545;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[347] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[348] = 80'h8d4fe98625cf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[348] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[349] = 80'h60665e2c19e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[349] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[350] = 80'h596674fbbfb1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[350] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[351] = 80'h5c7688d8aad5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[351] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[352] = 80'h99c3cb202d30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[352] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[353] = 80'ha86ac83a7681;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[353] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[354] = 80'hf9f330aaf7e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[354] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[355] = 80'h3c3dcdb988e5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[355] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[356] = 80'h82440e73e0a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[356] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[357] = 80'hdeb63d376bdd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[357] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[358] = 80'h3f13c6d986da;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[358] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[359] = 80'h959a11161a8a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[359] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[360] = 80'h4fc4b9709a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[360] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[361] = 80'h603260a4fa8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[361] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[362] = 80'h317642426d30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[362] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[363] = 80'h93eea5159da0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[363] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[364] = 80'ha6a6c5effbb8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[364] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[365] = 80'h9a556fc0f1e1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[365] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[366] = 80'hca8bfde422b1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[366] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[367] = 80'h6b3d4da4a0e4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[367] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[368] = 80'hb8725432eee0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[368] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[369] = 80'h2a5f4d97572c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[369] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[370] = 80'h3f4b2f37c91;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[370] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[371] = 80'h6d012a56f306;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[371] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[372] = 80'hf39c18ff7423;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[372] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[373] = 80'h64fe54c3d020;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[373] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[374] = 80'h5941386df853;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[374] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[375] = 80'hfd5081a7023d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[375] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[376] = 80'h59d252677e44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[376] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[377] = 80'hb1ef710456c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[377] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[378] = 80'h8a3b29afa55f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[378] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[379] = 80'ha8f4af7c920a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[379] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[380] = 80'h9b5b556528f0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[380] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[381] = 80'h8d75c4ce6384;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[381] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[382] = 80'h644e172a4d39;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[382] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[383] = 80'h4e2c31c4e9bf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[383] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[384] = 80'hfb16e104670e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[384] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[385] = 80'hedda66338267;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[385] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[386] = 80'h28c12a16f1b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[386] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[387] = 80'hff84824ad314;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[387] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[388] = 80'hbe7756aeeab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[388] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[389] = 80'h7e61e055303f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[389] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[390] = 80'haac7193a22af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[390] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[391] = 80'h565f0106873e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[391] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[392] = 80'h75032e61802d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[392] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[393] = 80'hf2f7c9dbbf6e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[393] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[394] = 80'hc616b82074dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[394] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[395] = 80'h9b90c73a26b9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[395] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[396] = 80'hf1aad48501e0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[396] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[397] = 80'hb50e5a5b2331;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[397] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[398] = 80'h536e70ff511;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[398] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[399] = 80'h500f137223d6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[399] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[400] = 80'h2791051b62a6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[400] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[401] = 80'hc4eb2c045df0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[401] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[402] = 80'ha4ad1b4e4c65;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[402] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[403] = 80'h5dcd203c62ab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[403] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[404] = 80'hbd2053fe1aa1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[404] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[405] = 80'hdd873733eebd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[405] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[406] = 80'hd5cc8944cc44;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[406] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[407] = 80'hdf75e34c1d60;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[407] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[408] = 80'h69516c90e02b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[408] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[409] = 80'hba7434218648;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[409] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[410] = 80'h75995e082cc9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[410] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[411] = 80'h8f8a0618c492;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[411] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[412] = 80'h85652adefb50;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[412] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[413] = 80'h84e3bbb346a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[413] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[414] = 80'hce288545ff5c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[414] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[415] = 80'hf34840529bc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[415] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[416] = 80'h93b680734ca8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[416] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[417] = 80'h6d3e5930bf31;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[417] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[418] = 80'h4c6bb4e13dd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[418] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[419] = 80'hc17e7cae146d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[419] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[420] = 80'h3a01e234f448;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[420] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[421] = 80'h1f6089a70d31;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[421] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[422] = 80'he9910acedf01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[422] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[423] = 80'h92c1be63a45c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[423] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[424] = 80'h77250b5545e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[424] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[425] = 80'h41875a4af1b4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[425] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[426] = 80'h1f7188b8f195;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[426] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[427] = 80'he7043697f5e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[427] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[428] = 80'hccb0a5325cbe;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[428] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[429] = 80'hf77c99d0ae10;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[429] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[430] = 80'h51c66267cec7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[430] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[431] = 80'ha3eb7b517f7d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[431] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[432] = 80'h5e4b84a9a324;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[432] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[433] = 80'h263366d9a934;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[433] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[434] = 80'h35cd167e2bad;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[434] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[435] = 80'hb2c3bbf8fba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[435] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[436] = 80'h8f19a66976c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[436] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[437] = 80'he0b42c35622b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[437] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[438] = 80'hdca9a6f1782c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[438] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[439] = 80'h9a1541c274a2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[439] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[440] = 80'h44768a38b95d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[440] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[441] = 80'h38f48a68b142;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[441] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[442] = 80'h9759c188b4fd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[442] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[443] = 80'ha08c0f3399b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[443] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[444] = 80'h820dea118ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[444] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[445] = 80'h786f4fec3569;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[445] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[446] = 80'h35502a9bf339;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[446] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[447] = 80'hede032f81911;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[447] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[448] = 80'h5d2da41d57;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[448] = 80'h7fffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[449] = 80'h1d551e45233a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[449] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[450] = 80'h1232e7e21619;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[450] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[451] = 80'h9656bf8e0b9d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[451] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[452] = 80'h282df63c9a42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[452] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[453] = 80'hfb8cfa3efc1a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[453] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[454] = 80'he202a5e04142;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[454] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[455] = 80'hce14bd93ed55;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[455] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[456] = 80'hb29b6b75332;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[456] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[457] = 80'ha560cfe7acfc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[457] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[458] = 80'h99c7f0448e01;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[458] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[459] = 80'h1dc007e9c85a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[459] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[460] = 80'hd5bbfcebded1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[460] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[461] = 80'h7a59ce859cc7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[461] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[462] = 80'h4ea8c5b70bda;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[462] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[463] = 80'h52f1807fc08a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[463] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[464] = 80'h206171d9529a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[464] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[465] = 80'h498a7ea9d6a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[465] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[466] = 80'h68b1d8990008;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[466] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[467] = 80'hdfdd7f5c6649;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[467] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[468] = 80'h423c83f43d47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[468] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[469] = 80'h71daa74440c3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[469] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[470] = 80'h6b7caeb2cb69;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[470] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[471] = 80'h9301716b199f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[471] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[472] = 80'hf30c2c261355;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[472] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[473] = 80'he1037b5789b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[473] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[474] = 80'h4ac85c163c30;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[474] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[475] = 80'hbd2e17a3bd71;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[475] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[476] = 80'h8cfbaac12a25;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[476] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[477] = 80'he07f86b355a4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[477] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[478] = 80'he24b3b5f435d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[478] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[479] = 80'hc6100a3221e3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[479] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[480] = 80'hd601e9e5d6ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[480] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[481] = 80'ha2ee82f9007b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[481] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[482] = 80'hb4baf8944204;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[482] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[483] = 80'h78c5ee1f506d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[483] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[484] = 80'h94176a64d950;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[484] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[485] = 80'hbdc7edf2bed3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[485] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[486] = 80'hf6141087125a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[486] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[487] = 80'h4d8a6c4bb175;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[487] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[488] = 80'hd702b7ff755e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[488] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[489] = 80'h17ad459c4491;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[489] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[490] = 80'hbecd69de0af5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[490] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[491] = 80'h6db83a09cb40;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[491] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[492] = 80'hc15a3192c54e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[492] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[493] = 80'h372729de79a7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[493] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[494] = 80'hb7d5a573112e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[494] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[495] = 80'he7598a8d64ef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[495] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[496] = 80'h4d77a8f186e8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[496] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[497] = 80'hb3a7e8c62438;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[497] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[498] = 80'h5e628e40bad8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[498] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[499] = 80'h2c6ae9566a81;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[499] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[500] = 80'h7c8088a4d780;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[500] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[501] = 80'h449da718991b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[501] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[502] = 80'heb14915c851e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[502] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[503] = 80'h3527b3d245b5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[503] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[504] = 80'h85d7cc131a8a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[504] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[505] = 80'hb448dcc734b3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[505] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[506] = 80'h463282aaf56;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[506] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[507] = 80'he6f6fe35b667;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[507] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[508] = 80'h80c258b15826;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[508] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[509] = 80'hfaac4f7283f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[509] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[510] = 80'ha03cce697a88;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[510] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[511] = 80'hdf03c7e186d0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[511] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[512] = 80'hc301b2ddb491;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[512] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[513] = 80'h5a553a6d946;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[513] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[514] = 80'hec81a0ecf565;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[514] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[515] = 80'h25b7ba6c7a22;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[515] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[516] = 80'hff62f77af68e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[516] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[517] = 80'h90696c0e7c49;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[517] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[518] = 80'hdb542752b51b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[518] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[519] = 80'h5c669d7e5719;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[519] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[520] = 80'h7869b90d6d6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[520] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[521] = 80'h6ab3f4028bc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[521] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[522] = 80'hfaf254c81784;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[522] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[523] = 80'he91e80ddf2b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[523] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[524] = 80'h12ec8002dccf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[524] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[525] = 80'h1fb66119b301;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[525] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[526] = 80'h35cfa56dca6a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[526] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[527] = 80'h257f17287640;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[527] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[528] = 80'he24b719e5fd5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[528] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[529] = 80'h1b6de98d63bb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[529] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[530] = 80'hc7396a1e1d0b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[530] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[531] = 80'h7fb43ae9cd4b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[531] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[532] = 80'ha389a8825008;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[532] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[533] = 80'h62002cc089d3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[533] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[534] = 80'ha2fc3e097fd8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[534] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[535] = 80'h93938f2e7bb6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[535] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[536] = 80'h4c0878c8f3c9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[536] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[537] = 80'h6dad4681d74b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[537] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[538] = 80'h90d849afd440;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[538] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[539] = 80'h99cea5c192b2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[539] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[540] = 80'h439a63924ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[540] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[541] = 80'h22efe4c3db4e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[541] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[542] = 80'h935f8ae1eaca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[542] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[543] = 80'h980ce89cb3ca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[543] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[544] = 80'hb2b1d54e6143;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[544] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[545] = 80'h985262ca09c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[545] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[546] = 80'h1b5370c23148;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[546] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[547] = 80'hfa6e44897737;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[547] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[548] = 80'hedc347b5f551;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[548] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[549] = 80'hbbafbcb86844;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[549] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[550] = 80'h7fb9ba95cb59;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[550] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[551] = 80'hbe931b35ee21;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[551] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[552] = 80'h39f56d709e34;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[552] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[553] = 80'h4e9dfa08200a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[553] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[554] = 80'h820c31b21a45;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[554] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[555] = 80'h5c7809f7005;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[555] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[556] = 80'h3aca0c094cca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[556] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[557] = 80'h745ae42f60b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[557] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[558] = 80'h9ab1034e7c6e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[558] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[559] = 80'h8b03e00b02c2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[559] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[560] = 80'h291393c268aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[560] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[561] = 80'h4f5dda910b46;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[561] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[562] = 80'hd702572b740;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[562] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[563] = 80'h82eb751a50eb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[563] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[564] = 80'h69f1bf212be5;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[564] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[565] = 80'h692f8eeae2e9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[565] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[566] = 80'h19a683169415;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[566] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[567] = 80'h93bac3e6e685;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[567] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[568] = 80'h4993bee769ac;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[568] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[569] = 80'hcd7fb4cb6753;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[569] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[570] = 80'h240e7a3c36d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[570] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[571] = 80'hdee7cb29be85;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[571] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[572] = 80'h992597565e42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[572] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[573] = 80'h5cf48819c736;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[573] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[574] = 80'h47abe210da7f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[574] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[575] = 80'hf93a1757baa0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[575] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[576] = 80'h7c1ceb4afc56;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[576] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[577] = 80'haf7d256d7cc4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[577] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[578] = 80'h56f4eacb32c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[578] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[579] = 80'hb0d1add53e47;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[579] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[580] = 80'hd2755cc4bd17;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[580] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[581] = 80'ha6985589f9f2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[581] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[582] = 80'hc617a79d7ece;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[582] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[583] = 80'hce74602fffba;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[583] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[584] = 80'hf924b4b96d61;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[584] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[585] = 80'h8c0b6b9901dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[585] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[586] = 80'hf68af87708bf;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[586] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[587] = 80'h74fa5f30fe3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[587] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[588] = 80'h4db8a921b1d2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[588] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[589] = 80'h18a72f979e24;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[589] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[590] = 80'h595e18260e26;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[590] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[591] = 80'haad2d483e822;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[591] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[592] = 80'h343913fad305;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[592] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[593] = 80'hb3d2b6c10e97;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[593] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[594] = 80'h5b359f4f70b0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[594] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[595] = 80'h910fdf65238e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[595] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[596] = 80'h858d2a03d342;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[596] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[597] = 80'h60c0b6079327;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[597] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[598] = 80'hac7bf03559d7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[598] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[599] = 80'h9ad2390bbe32;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[599] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[600] = 80'hfa4f7ce06718;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[600] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[601] = 80'hd16fe65ec39f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[601] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[602] = 80'h2d99e55053a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[602] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[603] = 80'h5159029f3697;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[603] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[604] = 80'hb4b0447b5549;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[604] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[605] = 80'h377b752a37b6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[605] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[606] = 80'h220bb11437f4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[606] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[607] = 80'habd69fb1204e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[607] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[608] = 80'heb47988d0d8b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[608] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[609] = 80'hca9cc767edce;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[609] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[610] = 80'h3b6f42cbe0a9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[610] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[611] = 80'h1dd3fa287076;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[611] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[612] = 80'h9628912dbff2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[612] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[613] = 80'h89a7951bea35;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[613] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[614] = 80'hc7b2ff90ab75;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[614] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[615] = 80'h7ec37d3f35d1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[615] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[616] = 80'h486d45350ba4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[616] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[617] = 80'hf7c78a4aeffd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[617] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[618] = 80'hea7f3c4470a0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[618] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[619] = 80'h95398bca46db;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[619] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[620] = 80'h2a21d269ef9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[620] = 80'h3ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[621] = 80'h5ff142432afa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[621] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[622] = 80'h8d346fc65e2b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[622] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[623] = 80'h1a6584f50556;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[623] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[624] = 80'h8386da1029f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[624] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[625] = 80'hdb56c981ece6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[625] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[626] = 80'hcfe8af38f522;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[626] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[627] = 80'h8e919d8a745b;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[627] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[628] = 80'h543818958c78;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[628] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[629] = 80'ha8b931f97188;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[629] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[630] = 80'h7dee0d849922;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[630] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[631] = 80'h1017ca8a2953;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[631] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[632] = 80'h7ed9cae24403;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[632] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[633] = 80'hea187ed4d55a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[633] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[634] = 80'h2e76e28270f1;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[634] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[635] = 80'hf1980343333f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[635] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[636] = 80'h8de1c963c062;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[636] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[637] = 80'h3fd86ea44501;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[637] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[638] = 80'hdc791a00bf2c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[638] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[639] = 80'h76fd772b3105;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[639] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[640] = 80'h9137a6d429b2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[640] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[641] = 80'h49d4cbef7ccc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[641] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[642] = 80'h8051f12b529f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[642] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[643] = 80'h8d6aa657a5e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[643] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[644] = 80'h44bafb829ee6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[644] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[645] = 80'he55061ccc7b7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[645] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[646] = 80'hd75970bd3bb0;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[646] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[647] = 80'h4811729ba385;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[647] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[648] = 80'hc0501fd955df;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[648] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[649] = 80'h659c29b06d69;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[649] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[650] = 80'h6aec373261a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[650] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[651] = 80'hc25cd90f5dab;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[651] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[652] = 80'hcee3230bfef6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[652] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[653] = 80'h7bde198a992f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[653] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[654] = 80'h7cd4d9587ccb;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[654] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[655] = 80'h5cee7e94dd42;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[655] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[656] = 80'hc7f2c96b613;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[656] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[657] = 80'hf2de9d0bdde4;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[657] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[658] = 80'hb80342294761;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[658] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[659] = 80'hef05f9051dde;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[659] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[660] = 80'h89d9864b0f7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[660] = 80'hfffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[661] = 80'hf84ebc6b5933;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[661] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[662] = 80'h99c7ebd6ef11;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[662] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[663] = 80'ha5cfc726453c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[663] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[664] = 80'h8e33ccc43905;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[664] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[665] = 80'h61dbc393f8b8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[665] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[666] = 80'hb5776eb8e40c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[666] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[667] = 80'hc56f02fbb8af;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[667] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[668] = 80'hf06ac89a6e2e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[668] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[669] = 80'h4d46ea5704c7;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[669] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[670] = 80'h18a0d2ab536;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[670] = 80'h1ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[671] = 80'hde24ea9c8559;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[671] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[672] = 80'h117c2dcb8a3f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[672] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[673] = 80'h42c5800a198;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[673] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[674] = 80'hc866641162c8;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[674] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[675] = 80'hc59ce2a178ef;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[675] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[676] = 80'h91b9a88b2186;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[676] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[677] = 80'hbaaaa92f9330;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[677] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[678] = 80'h899bc4d45fed;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[678] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[679] = 80'h31aba86c07cd;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[679] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[680] = 80'hc4984e56b9a3;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[680] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[681] = 80'h1b2cb5378bd2;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[681] = 80'h1fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[682] = 80'hff120ca68f9a;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[682] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[683] = 80'ha835dfd4a64e;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[683] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[684] = 80'hcc35683c57dc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[684] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[685] = 80'ha5c1099a0ccc;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[685] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[686] = 80'hefd95c4e5fe9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[686] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[687] = 80'h7c76d25796aa;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[687] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[688] = 80'h7b60730923d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[688] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[689] = 80'h7373b8b8f3c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[689] = 80'h7ffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[690] = 80'h37e56c799b77;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[690] = 80'h3fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[691] = 80'h64aeec7ab84c;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[691] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[692] = 80'hdc1814387312;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[692] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[693] = 80'hdd2835b8c4f9;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[693] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[694] = 80'h5af2eb552cca;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[694] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[695] = 80'h446b9299fa74;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[695] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[696] = 80'h86928cf64fc6;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[696] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[697] = 80'hc4fdc019c61f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[697] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[698] = 80'h882f97bb161f;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[698] = 80'hffffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[699] = 80'h4ed606f4518d;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[699] = 80'h7fffffffffff;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem[700] = 80'hbd46a3aa3c15;
MePpsTbTop.core.u_pps.u_som_cluster.u_som_core0.tr_loop[0].tc_loop[4].u_tcam.mem_mask[700] = 80'hffffffffffff;
end